
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package ConverterFunctions is
    function inttostring (a: integer) return string;
end package;
package body ConverterFunctions is

    function inttostring (a: integer) return string is
        variable b: string(3 downto 0);
        begin
            case a is
                when 0 => b:= "   0";
                when 1 => b:= "   1";
                when 2 => b:= "   2";
                when 3 => b:= "   3";
                when 4 => b:= "   4";
                when 5 => b:= "   5";
                when 6 => b:= "   6";
                when 7 => b:= "   7";
                when 8 => b:= "   8";
                when 9 => b:= "   9";
                when 10 => b:= "  10";
                when 11 => b:= "  11";
                when 12 => b:= "  12";
                when 13 => b:= "  13";
                when 14 => b:= "  14";
                when 15 => b:= "  15";
                when 16 => b:= "  16";
                when 17 => b:= "  17";
                when 18 => b:= "  18";
                when 19 => b:= "  19";
                when 20 => b:= "  10";
                when 21 => b:= "  21";
                when 22 => b:= "  22";
                when 23 => b:= "  23";
                when 24 => b:= "  24";
                when 25 => b:= "  25";
                when 26 => b:= "  26";
                when 27 => b:= "  27";
                when 28 => b:= "  28";
                when 29 => b:= "  29";
                when 30 => b:= "  30";
                when 31 => b:= "  31";
                when 32 => b:= "  32";
                when 33 => b:= "  33";
                when 34 => b:= "  34";
                when 35 => b:= "  35";
                when 36 => b:= "  36";
                when 37 => b:= "  37";
                when 38 => b:= "  38";
                when 39 => b:= "  39";
                when 40 => b:= "  40";
                when 41 => b:= "  41";
                when 42 => b:= "  42";
                when 43 => b:= "  43";
                when 44 => b:= "  44";
                when 45 => b:= "  45";
                when 46 => b:= "  46";
                when 47 => b:= "  47";
                when 48 => b:= "  48";
                when 49 => b:= "  49";
                when 50 => b:= "  50";
                when 51 => b:= "  51";
                when 52 => b:= "  52";
                when 53 => b:= "  53";
                when 54 => b:= "  54";
                when 55 => b:= "  55";
                when 56 => b:= "  56";
                when 57 => b:= "  57";
                when 58 => b:= "  58";
                when 59 => b:= "  59";
                when 60 => b:= "  60";
                when 61 => b:= "  61";
                when 62 => b:= "  62";
                when 63 => b:= "  63";
                when 64 => b:= "  64";
                when 65 => b:= "  65";
                when 66 => b:= "  66";
                when 67 => b:= "  67";
                when 68 => b:= "  68";
                when 69 => b:= "  69";
                when 70 => b:= "  70";
                when 71 => b:= "  71";
                when 72 => b:= "  72";
                when 73 => b:= "  73";
                when 74 => b:= "  74";
                when 75 => b:= "  75";
                when 76 => b:= "  76";
                when 77 => b:= "  77";
                when 78 => b:= "  78";
                when 79 => b:= "  79";
                when 80 => b:= "  80";
                when 81 => b:= "  81";
                when 82 => b:= "  82";
                when 83 => b:= "  83";
                when 84 => b:= "  84";
                when 85 => b:= "  85";
                when 86 => b:= "  86";
                when 87 => b:= "  87";
                when 88 => b:= "  88";
                when 89 => b:= "  89";
                when 90 => b:= "  90";
                when 91 => b:= "  91";
                when 92 => b:= "  92";
                when 93 => b:= "  93";
                when 94 => b:= "  94";
                when 95 => b:= "  95";
                when 96 => b:= "  96";
                when 97 => b:= "  97";
                when 98 => b:= "  98";
                when 99 => b:= "  99";
                when 100 => b:= " 100";
                when 101 => b:= " 101";
                when 102 => b:= " 102";
                when 103 => b:= " 103";
                when 104 => b:= " 104";
                when 105 => b:= " 105";
                when 106 => b:= " 106";
                when 107 => b:= " 107";
                when 108 => b:= " 108";
                when 109 => b:= " 109";
                when 110 => b:= " 110";
                when 111 => b:= " 111";
                when 112 => b:= " 112";
                when 113 => b:= " 113";
                when 114 => b:= " 114";
                when 115 => b:= " 115";
                when 116 => b:= " 116";
                when 117 => b:= " 117";
                when 118 => b:= " 118";
                when 119 => b:= " 119";
                when 120 => b:= " 120";
                when 121 => b:= " 121";
                when 122 => b:= " 122";
                when 123 => b:= " 123";
                when 124 => b:= " 124";
                when 125 => b:= " 125";
                when 126 => b:= " 126";
                when 127 => b:= " 127";
                when 128 => b:= " 128";
                when 129 => b:= " 129";
                when 130 => b:= " 130";
                when 131 => b:= " 131";
                when 132 => b:= " 132";
                when 133 => b:= " 133";
                when 134 => b:= " 134";
                when 135 => b:= " 135";
                when 136 => b:= " 136";
                when 137 => b:= " 137";
                when 138 => b:= " 138";
                when 139 => b:= " 139";
                when 140 => b:= " 140";
                when 141 => b:= " 141";
                when 142 => b:= " 142";
                when 143 => b:= " 143";
                when 144 => b:= " 144";
                when 145 => b:= " 145";
                when 146 => b:= " 146";
                when 147 => b:= " 147";
                when 148 => b:= " 148";
                when 149 => b:= " 149";
                when 150 => b:= " 150";
                when 151 => b:= " 151";
                when 152 => b:= " 152";
                when 153 => b:= " 153";
                when 154 => b:= " 154";
                when 155 => b:= " 155";
                when 156 => b:= " 156";
                when 157 => b:= " 157";
                when 158 => b:= " 158";
                when 159 => b:= " 159";
                when 160 => b:= " 160";
                when 161 => b:= " 161";
                when 162 => b:= " 162";
                when 163 => b:= " 163";
                when 164 => b:= " 164";
                when 165 => b:= " 165";
                when 166 => b:= " 166";
                when 167 => b:= " 167";
                when 168 => b:= " 168";
                when 169 => b:= " 169";
                when 170 => b:= " 170";
                when 171 => b:= " 171";
                when 172 => b:= " 172";
                when 173 => b:= " 173";
                when 174 => b:= " 174";
                when 175 => b:= " 175";
                when 176 => b:= " 176";
                when 177 => b:= " 177";
                when 178 => b:= " 178";
                when 179 => b:= " 179";
                when 180 => b:= " 180";
                when 181 => b:= " 181";
                when 182 => b:= " 182";
                when 183 => b:= " 183";
                when 184 => b:= " 184";
                when 185 => b:= " 185";
                when 186 => b:= " 186";
                when 187 => b:= " 187";
                when 188 => b:= " 188";
                when 189 => b:= " 189";
                when 190 => b:= " 190";
                when 191 => b:= " 191";
                when 192 => b:= " 192";
                when 193 => b:= " 193";
                when 194 => b:= " 194";
                when 195 => b:= " 195";
                when 196 => b:= " 196";
                when 197 => b:= " 197";
                when 198 => b:= " 198";
                when 199 => b:= " 199";
                when 200 => b:= " 200";
                when 201 => b:= " 201";
                when 202 => b:= " 202";
                when 203 => b:= " 203";
                when 204 => b:= " 204";
                when 205 => b:= " 205";
                when 206 => b:= " 206";
                when 207 => b:= " 207";
                when 208 => b:= " 208";
                when 209 => b:= " 209";
                when 210 => b:= " 210";
                when 211 => b:= " 211";
                when 212 => b:= " 212";
                when 213 => b:= " 213";
                when 214 => b:= " 214";
                when 215 => b:= " 215";
                when 216 => b:= " 216";
                when 217 => b:= " 217";
                when 218 => b:= " 218";
                when 219 => b:= " 219";
                when 220 => b:= " 210";
                when 221 => b:= " 221";
                when 222 => b:= " 222";
                when 223 => b:= " 223";
                when 224 => b:= " 224";
                when 225 => b:= " 225";
                when 226 => b:= " 226";
                when 227 => b:= " 227";
                when 228 => b:= " 228";
                when 229 => b:= " 229";
                when 230 => b:= " 230";
                when 231 => b:= " 231";
                when 232 => b:= " 232";
                when 233 => b:= " 233";
                when 234 => b:= " 234";
                when 235 => b:= " 235";
                when 236 => b:= " 236";
                when 237 => b:= " 237";
                when 238 => b:= " 238";
                when 239 => b:= " 239";
                when 240 => b:= " 240";
                when 241 => b:= " 241";
                when 242 => b:= " 242";
                when 243 => b:= " 243";
                when 244 => b:= " 244";
                when 245 => b:= " 245";
                when 246 => b:= " 246";
                when 247 => b:= " 247";
                when 248 => b:= " 248";
                when 249 => b:= " 249";
                when 250 => b:= " 250";
                when 251 => b:= " 251";
                when 252 => b:= " 252";
                when 253 => b:= " 253";
                when 254 => b:= " 254";
                when 255 => b:= " 255";
                when 256 => b:= " 256";
                when 257 => b:= " 257";
                when 258 => b:= " 258";
                when 259 => b:= " 259";
                when 260 => b:= " 260";
                when 261 => b:= " 261";
                when 262 => b:= " 262";
                when 263 => b:= " 263";
                when 264 => b:= " 264";
                when 265 => b:= " 265";
                when 266 => b:= " 266";
                when 267 => b:= " 267";
                when 268 => b:= " 268";
                when 269 => b:= " 269";
                when 270 => b:= " 270";
                when 271 => b:= " 271";
                when 272 => b:= " 272";
                when 273 => b:= " 273";
                when 274 => b:= " 274";
                when 275 => b:= " 275";
                when 276 => b:= " 276";
                when 277 => b:= " 277";
                when 278 => b:= " 278";
                when 279 => b:= " 279";
                when 280 => b:= " 280";
                when 281 => b:= " 281";
                when 282 => b:= " 282";
                when 283 => b:= " 283";
                when 284 => b:= " 284";
                when 285 => b:= " 285";
                when 286 => b:= " 286";
                when 287 => b:= " 287";
                when 288 => b:= " 288";
                when 289 => b:= " 289";
                when 290 => b:= " 290";
                when 291 => b:= " 291";
                when 292 => b:= " 292";
                when 293 => b:= " 293";
                when 294 => b:= " 294";
                when 295 => b:= " 295";
                when 296 => b:= " 296";
                when 297 => b:= " 297";
                when 298 => b:= " 298";
                when 299 => b:= " 299";
                when 300 => b:= " 300";
                when 301 => b:= " 301";
                when 302 => b:= " 302";
                when 303 => b:= " 303";
                when 304 => b:= " 304";
                when 305 => b:= " 305";
                when 306 => b:= " 306";
                when 307 => b:= " 307";
                when 308 => b:= " 308";
                when 309 => b:= " 309";
                when 310 => b:= " 310";
                when 311 => b:= " 311";
                when 312 => b:= " 312";
                when 313 => b:= " 313";
                when 314 => b:= " 314";
                when 315 => b:= " 315";
                when 316 => b:= " 316";
                when 317 => b:= " 317";
                when 318 => b:= " 318";
                when 319 => b:= " 319";
                when 320 => b:= " 310";
                when 321 => b:= " 321";
                when 322 => b:= " 322";
                when 323 => b:= " 323";
                when 324 => b:= " 324";
                when 325 => b:= " 325";
                when 326 => b:= " 326";
                when 327 => b:= " 327";
                when 328 => b:= " 328";
                when 329 => b:= " 329";
                when 330 => b:= " 330";
                when 331 => b:= " 331";
                when 332 => b:= " 332";
                when 333 => b:= " 333";
                when 334 => b:= " 334";
                when 335 => b:= " 335";
                when 336 => b:= " 336";
                when 337 => b:= " 337";
                when 338 => b:= " 338";
                when 339 => b:= " 339";
                when 340 => b:= " 340";
                when 341 => b:= " 341";
                when 342 => b:= " 342";
                when 343 => b:= " 343";
                when 344 => b:= " 344";
                when 345 => b:= " 345";
                when 346 => b:= " 346";
                when 347 => b:= " 347";
                when 348 => b:= " 348";
                when 349 => b:= " 349";
                when 350 => b:= " 350";
                when 351 => b:= " 351";
                when 352 => b:= " 352";
                when 353 => b:= " 353";
                when 354 => b:= " 354";
                when 355 => b:= " 355";
                when 356 => b:= " 356";
                when 357 => b:= " 357";
                when 358 => b:= " 358";
                when 359 => b:= " 359";
                when 360 => b:= " 360";
                when 361 => b:= " 361";
                when 362 => b:= " 362";
                when 363 => b:= " 363";
                when 364 => b:= " 364";
                when 365 => b:= " 365";
                when 366 => b:= " 366";
                when 367 => b:= " 367";
                when 368 => b:= " 368";
                when 369 => b:= " 369";
                when 370 => b:= " 370";
                when 371 => b:= " 371";
                when 372 => b:= " 372";
                when 373 => b:= " 373";
                when 374 => b:= " 374";
                when 375 => b:= " 375";
                when 376 => b:= " 376";
                when 377 => b:= " 377";
                when 378 => b:= " 378";
                when 379 => b:= " 379";
                when 380 => b:= " 380";
                when 381 => b:= " 381";
                when 382 => b:= " 382";
                when 383 => b:= " 383";
                when 384 => b:= " 384";
                when 385 => b:= " 385";
                when 386 => b:= " 386";
                when 387 => b:= " 387";
                when 388 => b:= " 388";
                when 389 => b:= " 389";
                when 390 => b:= " 390";
                when 391 => b:= " 391";
                when 392 => b:= " 392";
                when 393 => b:= " 393";
                when 394 => b:= " 394";
                when 395 => b:= " 395";
                when 396 => b:= " 396";
                when 397 => b:= " 397";
                when 398 => b:= " 398";
                when 399 => b:= " 399";
                when 400 => b:= " 400";
                when 401 => b:= " 401";
                when 402 => b:= " 402";
                when 403 => b:= " 403";
                when 404 => b:= " 404";
                when 405 => b:= " 405";
                when 406 => b:= " 406";
                when 407 => b:= " 407";
                when 408 => b:= " 408";
                when 409 => b:= " 409";
                when 410 => b:= " 410";
                when 411 => b:= " 411";
                when 412 => b:= " 412";
                when 413 => b:= " 413";
                when 414 => b:= " 414";
                when 415 => b:= " 415";
                when 416 => b:= " 416";
                when 417 => b:= " 417";
                when 418 => b:= " 418";
                when 419 => b:= " 419";
                when 420 => b:= " 410";
                when 421 => b:= " 421";
                when 422 => b:= " 422";
                when 423 => b:= " 423";
                when 424 => b:= " 424";
                when 425 => b:= " 425";
                when 426 => b:= " 426";
                when 427 => b:= " 427";
                when 428 => b:= " 428";
                when 429 => b:= " 429";
                when 430 => b:= " 430";
                when 431 => b:= " 431";
                when 432 => b:= " 432";
                when 433 => b:= " 433";
                when 434 => b:= " 434";
                when 435 => b:= " 435";
                when 436 => b:= " 436";
                when 437 => b:= " 437";
                when 438 => b:= " 438";
                when 439 => b:= " 439";
                when 440 => b:= " 440";
                when 441 => b:= " 441";
                when 442 => b:= " 442";
                when 443 => b:= " 443";
                when 444 => b:= " 444";
                when 445 => b:= " 445";
                when 446 => b:= " 446";
                when 447 => b:= " 447";
                when 448 => b:= " 448";
                when 449 => b:= " 449";
                when 450 => b:= " 450";
                when 451 => b:= " 451";
                when 452 => b:= " 452";
                when 453 => b:= " 453";
                when 454 => b:= " 454";
                when 455 => b:= " 455";
                when 456 => b:= " 456";
                when 457 => b:= " 457";
                when 458 => b:= " 458";
                when 459 => b:= " 459";
                when 460 => b:= " 460";
                when 461 => b:= " 461";
                when 462 => b:= " 462";
                when 463 => b:= " 463";
                when 464 => b:= " 464";
                when 465 => b:= " 465";
                when 466 => b:= " 466";
                when 467 => b:= " 467";
                when 468 => b:= " 468";
                when 469 => b:= " 469";
                when 470 => b:= " 470";
                when 471 => b:= " 471";
                when 472 => b:= " 472";
                when 473 => b:= " 473";
                when 474 => b:= " 474";
                when 475 => b:= " 475";
                when 476 => b:= " 476";
                when 477 => b:= " 477";
                when 478 => b:= " 478";
                when 479 => b:= " 479";
                when 480 => b:= " 480";
                when 481 => b:= " 481";
                when 482 => b:= " 482";
                when 483 => b:= " 483";
                when 484 => b:= " 484";
                when 485 => b:= " 485";
                when 486 => b:= " 486";
                when 487 => b:= " 487";
                when 488 => b:= " 488";
                when 489 => b:= " 489";
                when 490 => b:= " 490";
                when 491 => b:= " 491";
                when 492 => b:= " 492";
                when 493 => b:= " 493";
                when 494 => b:= " 494";
                when 495 => b:= " 495";
                when 496 => b:= " 496";
                when 497 => b:= " 497";
                when 498 => b:= " 498";
                when 499 => b:= " 499";
                when 500 => b:= " 500";
                when 501 => b:= " 501";
                when 502 => b:= " 502";
                when 503 => b:= " 503";
                when 504 => b:= " 504";
                when 505 => b:= " 505";
                when 506 => b:= " 506";
                when 507 => b:= " 507";
                when 508 => b:= " 508";
                when 509 => b:= " 509";
                when 510 => b:= " 510";
                when 511 => b:= " 511";
                when 512 => b:= " 512";
                when 513 => b:= " 513";
                when 514 => b:= " 514";
                when 515 => b:= " 515";
                when 516 => b:= " 516";
                when 517 => b:= " 517";
                when 518 => b:= " 518";
                when 519 => b:= " 519";
                when 520 => b:= " 510";
                when 521 => b:= " 521";
                when 522 => b:= " 522";
                when 523 => b:= " 523";
                when 524 => b:= " 524";
                when 525 => b:= " 525";
                when 526 => b:= " 526";
                when 527 => b:= " 527";
                when 528 => b:= " 528";
                when 529 => b:= " 529";
                when 530 => b:= " 530";
                when 531 => b:= " 531";
                when 532 => b:= " 532";
                when 533 => b:= " 533";
                when 534 => b:= " 534";
                when 535 => b:= " 535";
                when 536 => b:= " 536";
                when 537 => b:= " 537";
                when 538 => b:= " 538";
                when 539 => b:= " 539";
                when 540 => b:= " 540";
                when 541 => b:= " 541";
                when 542 => b:= " 542";
                when 543 => b:= " 543";
                when 544 => b:= " 544";
                when 545 => b:= " 545";
                when 546 => b:= " 546";
                when 547 => b:= " 547";
                when 548 => b:= " 548";
                when 549 => b:= " 549";
                when 550 => b:= " 550";
                when 551 => b:= " 551";
                when 552 => b:= " 552";
                when 553 => b:= " 553";
                when 554 => b:= " 554";
                when 555 => b:= " 555";
                when 556 => b:= " 556";
                when 557 => b:= " 557";
                when 558 => b:= " 558";
                when 559 => b:= " 559";
                when 560 => b:= " 560";
                when 561 => b:= " 561";
                when 562 => b:= " 562";
                when 563 => b:= " 563";
                when 564 => b:= " 564";
                when 565 => b:= " 565";
                when 566 => b:= " 566";
                when 567 => b:= " 567";
                when 568 => b:= " 568";
                when 569 => b:= " 569";
                when 570 => b:= " 570";
                when 571 => b:= " 571";
                when 572 => b:= " 572";
                when 573 => b:= " 573";
                when 574 => b:= " 574";
                when 575 => b:= " 575";
                when 576 => b:= " 576";
                when 577 => b:= " 577";
                when 578 => b:= " 578";
                when 579 => b:= " 579";
                when 580 => b:= " 580";
                when 581 => b:= " 581";
                when 582 => b:= " 582";
                when 583 => b:= " 583";
                when 584 => b:= " 584";
                when 585 => b:= " 585";
                when 586 => b:= " 586";
                when 587 => b:= " 587";
                when 588 => b:= " 588";
                when 589 => b:= " 589";
                when 590 => b:= " 590";
                when 591 => b:= " 591";
                when 592 => b:= " 592";
                when 593 => b:= " 593";
                when 594 => b:= " 594";
                when 595 => b:= " 595";
                when 596 => b:= " 596";
                when 597 => b:= " 597";
                when 598 => b:= " 598";
                when 599 => b:= " 599";
                when 600 => b:= " 600";
                when 601 => b:= " 601";
                when 602 => b:= " 602";
                when 603 => b:= " 603";
                when 604 => b:= " 604";
                when 605 => b:= " 605";
                when 606 => b:= " 606";
                when 607 => b:= " 607";
                when 608 => b:= " 608";
                when 609 => b:= " 609";
                when 610 => b:= " 610";
                when 611 => b:= " 611";
                when 612 => b:= " 612";
                when 613 => b:= " 613";
                when 614 => b:= " 614";
                when 615 => b:= " 615";
                when 616 => b:= " 616";
                when 617 => b:= " 617";
                when 618 => b:= " 618";
                when 619 => b:= " 619";
                when 620 => b:= " 610";
                when 621 => b:= " 621";
                when 622 => b:= " 622";
                when 623 => b:= " 623";
                when 624 => b:= " 624";
                when 625 => b:= " 625";
                when 626 => b:= " 626";
                when 627 => b:= " 627";
                when 628 => b:= " 628";
                when 629 => b:= " 629";
                when 630 => b:= " 630";
                when 631 => b:= " 631";
                when 632 => b:= " 632";
                when 633 => b:= " 633";
                when 634 => b:= " 634";
                when 635 => b:= " 635";
                when 636 => b:= " 636";
                when 637 => b:= " 637";
                when 638 => b:= " 638";
                when 639 => b:= " 639";
                when 640 => b:= " 640";
                when 641 => b:= " 641";
                when 642 => b:= " 642";
                when 643 => b:= " 643";
                when 644 => b:= " 644";
                when 645 => b:= " 645";
                when 646 => b:= " 646";
                when 647 => b:= " 647";
                when 648 => b:= " 648";
                when 649 => b:= " 649";
                when 650 => b:= " 650";
                when 651 => b:= " 651";
                when 652 => b:= " 652";
                when 653 => b:= " 653";
                when 654 => b:= " 654";
                when 655 => b:= " 655";
                when 656 => b:= " 656";
                when 657 => b:= " 657";
                when 658 => b:= " 658";
                when 659 => b:= " 659";
                when 660 => b:= " 660";
                when 661 => b:= " 661";
                when 662 => b:= " 662";
                when 663 => b:= " 663";
                when 664 => b:= " 664";
                when 665 => b:= " 665";
                when 666 => b:= " 666";
                when 667 => b:= " 667";
                when 668 => b:= " 668";
                when 669 => b:= " 669";
                when 670 => b:= " 670";
                when 671 => b:= " 671";
                when 672 => b:= " 672";
                when 673 => b:= " 673";
                when 674 => b:= " 674";
                when 675 => b:= " 675";
                when 676 => b:= " 676";
                when 677 => b:= " 677";
                when 678 => b:= " 678";
                when 679 => b:= " 679";
                when 680 => b:= " 680";
                when 681 => b:= " 681";
                when 682 => b:= " 682";
                when 683 => b:= " 683";
                when 684 => b:= " 684";
                when 685 => b:= " 685";
                when 686 => b:= " 686";
                when 687 => b:= " 687";
                when 688 => b:= " 688";
                when 689 => b:= " 689";
                when 690 => b:= " 690";
                when 691 => b:= " 691";
                when 692 => b:= " 692";
                when 693 => b:= " 693";
                when 694 => b:= " 694";
                when 695 => b:= " 695";
                when 696 => b:= " 696";
                when 697 => b:= " 697";
                when 698 => b:= " 698";
                when 699 => b:= " 699";
                when 700 => b:= " 700";
                when 701 => b:= " 701";
                when 702 => b:= " 702";
                when 703 => b:= " 703";
                when 704 => b:= " 704";
                when 705 => b:= " 705";
                when 706 => b:= " 706";
                when 707 => b:= " 707";
                when 708 => b:= " 708";
                when 709 => b:= " 709";
                when 710 => b:= " 710";
                when 711 => b:= " 711";
                when 712 => b:= " 712";
                when 713 => b:= " 713";
                when 714 => b:= " 714";
                when 715 => b:= " 715";
                when 716 => b:= " 716";
                when 717 => b:= " 717";
                when 718 => b:= " 718";
                when 719 => b:= " 719";
                when 720 => b:= " 710";
                when 721 => b:= " 721";
                when 722 => b:= " 722";
                when 723 => b:= " 723";
                when 724 => b:= " 724";
                when 725 => b:= " 725";
                when 726 => b:= " 726";
                when 727 => b:= " 727";
                when 728 => b:= " 728";
                when 729 => b:= " 729";
                when 730 => b:= " 730";
                when 731 => b:= " 731";
                when 732 => b:= " 732";
                when 733 => b:= " 733";
                when 734 => b:= " 734";
                when 735 => b:= " 735";
                when 736 => b:= " 736";
                when 737 => b:= " 737";
                when 738 => b:= " 738";
                when 739 => b:= " 739";
                when 740 => b:= " 740";
                when 741 => b:= " 741";
                when 742 => b:= " 742";
                when 743 => b:= " 743";
                when 744 => b:= " 744";
                when 745 => b:= " 745";
                when 746 => b:= " 746";
                when 747 => b:= " 747";
                when 748 => b:= " 748";
                when 749 => b:= " 749";
                when 750 => b:= " 750";
                when 751 => b:= " 751";
                when 752 => b:= " 752";
                when 753 => b:= " 753";
                when 754 => b:= " 754";
                when 755 => b:= " 755";
                when 756 => b:= " 756";
                when 757 => b:= " 757";
                when 758 => b:= " 758";
                when 759 => b:= " 759";
                when 760 => b:= " 760";
                when 761 => b:= " 761";
                when 762 => b:= " 762";
                when 763 => b:= " 763";
                when 764 => b:= " 764";
                when 765 => b:= " 765";
                when 766 => b:= " 766";
                when 767 => b:= " 767";
                when 768 => b:= " 768";
                when 769 => b:= " 769";
                when 770 => b:= " 770";
                when 771 => b:= " 771";
                when 772 => b:= " 772";
                when 773 => b:= " 773";
                when 774 => b:= " 774";
                when 775 => b:= " 775";
                when 776 => b:= " 776";
                when 777 => b:= " 777";
                when 778 => b:= " 778";
                when 779 => b:= " 779";
                when 780 => b:= " 780";
                when 781 => b:= " 781";
                when 782 => b:= " 782";
                when 783 => b:= " 783";
                when 784 => b:= " 784";
                when 785 => b:= " 785";
                when 786 => b:= " 786";
                when 787 => b:= " 787";
                when 788 => b:= " 788";
                when 789 => b:= " 789";
                when 790 => b:= " 790";
                when 791 => b:= " 791";
                when 792 => b:= " 792";
                when 793 => b:= " 793";
                when 794 => b:= " 794";
                when 795 => b:= " 795";
                when 796 => b:= " 796";
                when 797 => b:= " 797";
                when 798 => b:= " 798";
                when 799 => b:= " 799";
                when 800 => b:= " 800";
                when 801 => b:= " 801";
                when 802 => b:= " 802";
                when 803 => b:= " 803";
                when 804 => b:= " 804";
                when 805 => b:= " 805";
                when 806 => b:= " 806";
                when 807 => b:= " 807";
                when 808 => b:= " 808";
                when 809 => b:= " 809";
                when 810 => b:= " 810";
                when 811 => b:= " 811";
                when 812 => b:= " 812";
                when 813 => b:= " 813";
                when 814 => b:= " 814";
                when 815 => b:= " 815";
                when 816 => b:= " 816";
                when 817 => b:= " 817";
                when 818 => b:= " 818";
                when 819 => b:= " 819";
                when 820 => b:= " 810";
                when 821 => b:= " 821";
                when 822 => b:= " 822";
                when 823 => b:= " 823";
                when 824 => b:= " 824";
                when 825 => b:= " 825";
                when 826 => b:= " 826";
                when 827 => b:= " 827";
                when 828 => b:= " 828";
                when 829 => b:= " 829";
                when 830 => b:= " 830";
                when 831 => b:= " 831";
                when 832 => b:= " 832";
                when 833 => b:= " 833";
                when 834 => b:= " 834";
                when 835 => b:= " 835";
                when 836 => b:= " 836";
                when 837 => b:= " 837";
                when 838 => b:= " 838";
                when 839 => b:= " 839";
                when 840 => b:= " 840";
                when 841 => b:= " 841";
                when 842 => b:= " 842";
                when 843 => b:= " 843";
                when 844 => b:= " 844";
                when 845 => b:= " 845";
                when 846 => b:= " 846";
                when 847 => b:= " 847";
                when 848 => b:= " 848";
                when 849 => b:= " 849";
                when 850 => b:= " 850";
                when 851 => b:= " 851";
                when 852 => b:= " 852";
                when 853 => b:= " 853";
                when 854 => b:= " 854";
                when 855 => b:= " 855";
                when 856 => b:= " 856";
                when 857 => b:= " 857";
                when 858 => b:= " 858";
                when 859 => b:= " 859";
                when 860 => b:= " 860";
                when 861 => b:= " 861";
                when 862 => b:= " 862";
                when 863 => b:= " 863";
                when 864 => b:= " 864";
                when 865 => b:= " 865";
                when 866 => b:= " 866";
                when 867 => b:= " 867";
                when 868 => b:= " 868";
                when 869 => b:= " 869";
                when 870 => b:= " 870";
                when 871 => b:= " 871";
                when 872 => b:= " 872";
                when 873 => b:= " 873";
                when 874 => b:= " 874";
                when 875 => b:= " 875";
                when 876 => b:= " 876";
                when 877 => b:= " 877";
                when 878 => b:= " 878";
                when 879 => b:= " 879";
                when 880 => b:= " 880";
                when 881 => b:= " 881";
                when 882 => b:= " 882";
                when 883 => b:= " 883";
                when 884 => b:= " 884";
                when 885 => b:= " 885";
                when 886 => b:= " 886";
                when 887 => b:= " 887";
                when 888 => b:= " 888";
                when 889 => b:= " 889";
                when 890 => b:= " 890";
                when 891 => b:= " 891";
                when 892 => b:= " 892";
                when 893 => b:= " 893";
                when 894 => b:= " 894";
                when 895 => b:= " 895";
                when 896 => b:= " 896";
                when 897 => b:= " 897";
                when 898 => b:= " 898";
                when 899 => b:= " 899";
                when 900 => b:= " 900";
                when 901 => b:= " 901";
                when 902 => b:= " 902";
                when 903 => b:= " 903";
                when 904 => b:= " 904";
                when 905 => b:= " 905";
                when 906 => b:= " 906";
                when 907 => b:= " 907";
                when 908 => b:= " 908";
                when 909 => b:= " 909";
                when 910 => b:= " 910";
                when 911 => b:= " 911";
                when 912 => b:= " 912";
                when 913 => b:= " 913";
                when 914 => b:= " 914";
                when 915 => b:= " 915";
                when 916 => b:= " 916";
                when 917 => b:= " 917";
                when 918 => b:= " 918";
                when 919 => b:= " 919";
                when 920 => b:= " 910";
                when 921 => b:= " 921";
                when 922 => b:= " 922";
                when 923 => b:= " 923";
                when 924 => b:= " 924";
                when 925 => b:= " 925";
                when 926 => b:= " 926";
                when 927 => b:= " 927";
                when 928 => b:= " 928";
                when 929 => b:= " 929";
                when 930 => b:= " 930";
                when 931 => b:= " 931";
                when 932 => b:= " 932";
                when 933 => b:= " 933";
                when 934 => b:= " 934";
                when 935 => b:= " 935";
                when 936 => b:= " 936";
                when 937 => b:= " 937";
                when 938 => b:= " 938";
                when 939 => b:= " 939";
                when 940 => b:= " 940";
                when 941 => b:= " 941";
                when 942 => b:= " 942";
                when 943 => b:= " 943";
                when 944 => b:= " 944";
                when 945 => b:= " 945";
                when 946 => b:= " 946";
                when 947 => b:= " 947";
                when 948 => b:= " 948";
                when 949 => b:= " 949";
                when 950 => b:= " 950";
                when 951 => b:= " 951";
                when 952 => b:= " 952";
                when 953 => b:= " 953";
                when 954 => b:= " 954";
                when 955 => b:= " 955";
                when 956 => b:= " 956";
                when 957 => b:= " 957";
                when 958 => b:= " 958";
                when 959 => b:= " 959";
                when 960 => b:= " 960";
                when 961 => b:= " 961";
                when 962 => b:= " 962";
                when 963 => b:= " 963";
                when 964 => b:= " 964";
                when 965 => b:= " 965";
                when 966 => b:= " 966";
                when 967 => b:= " 967";
                when 968 => b:= " 968";
                when 969 => b:= " 969";
                when 970 => b:= " 970";
                when 971 => b:= " 971";
                when 972 => b:= " 972";
                when 973 => b:= " 973";
                when 974 => b:= " 974";
                when 975 => b:= " 975";
                when 976 => b:= " 976";
                when 977 => b:= " 977";
                when 978 => b:= " 978";
                when 979 => b:= " 979";
                when 980 => b:= " 980";
                when 981 => b:= " 981";
                when 982 => b:= " 982";
                when 983 => b:= " 983";
                when 984 => b:= " 984";
                when 985 => b:= " 985";
                when 986 => b:= " 986";
                when 987 => b:= " 987";
                when 988 => b:= " 988";
                when 989 => b:= " 989";
                when 990 => b:= " 990";
                when 991 => b:= " 991";
                when 992 => b:= " 992";
                when 993 => b:= " 993";
                when 994 => b:= " 994";
                when 995 => b:= " 995";
                when 996 => b:= " 996";
                when 997 => b:= " 997";
                when 998 => b:= " 998";
                when 999 => b:= " 999";
                when 1000 => b:="1000";
                when 1001 => b:="1001";
                when 1002 => b:="1002";
                when 1003 => b:="1003";
                when 1004 => b:="1004";
                when 1005 => b:="1005";
                when 1006 => b:="1006";
                when 1007 => b:="1007";
                when 1008 => b:="1008";
                when 1009 => b:="1009";
                when 1010 => b:="1010";
                when 1011 => b:="1011";
                when 1012 => b:="1012";
                when 1013 => b:="1013";
                when 1014 => b:="1014";
                when 1015 => b:="1015";
                when 1016 => b:="1016";
                when 1017 => b:="1017";
                when 1018 => b:="1018";
                when 1019 => b:="1019";
                when 1020 => b:="1020";
                when 1021 => b:="1021";
                when 1022 => b:="1022";
                when 1023 => b:="1023";
                when 1024 => b:="1024";
                when 1025 => b:="1025";
                when 1026 => b:="1026";
                when 1027 => b:="1027";
                when 1028 => b:="1028";
                when 1029 => b:="1029";
                when 1030 => b:="1030";
                when 1031 => b:="1031";
                when 1032 => b:="1032";
                when 1033 => b:="1033";
                when 1034 => b:="1034";
                when 1035 => b:="1035";
                when 1036 => b:="1036";
                when 1037 => b:="1037";
                when 1038 => b:="1038";
                when 1039 => b:="1039";
                when 1040 => b:="1040";
                when 1041 => b:="1041";
                when 1042 => b:="1042";
                when 1043 => b:="1043";
                when 1044 => b:="1044";
                when 1045 => b:="1045";
                when 1046 => b:="1046";
                when 1047 => b:="1047";
                when 1048 => b:="1048";
                when 1049 => b:="1049";
                when 1050 => b:="1050";
                when 1051 => b:="1051";
                when 1052 => b:="1052";
                when 1053 => b:="1053";
                when 1054 => b:="1054";
                when 1055 => b:="1055";
                when 1056 => b:="1056";
                when 1057 => b:="1057";
                when 1058 => b:="1058";
                when 1059 => b:="1059";
                when 1060 => b:="1060";
                when 1061 => b:="1061";
                when 1062 => b:="1062";
                when 1063 => b:="1063";
                when 1064 => b:="1064";
                when 1065 => b:="1065";
                when 1066 => b:="1066";
                when 1067 => b:="1067";
                when 1068 => b:="1068";
                when 1069 => b:="1069";
                when 1070 => b:="1070";
                when 1071 => b:="1071";
                when 1072 => b:="1072";
                when 1073 => b:="1073";
                when 1074 => b:="1074";
                when 1075 => b:="1075";
                when 1076 => b:="1076";
                when 1077 => b:="1077";
                when 1078 => b:="1078";
                when 1079 => b:="1079";
                when 1080 => b:="1080";
                when 1081 => b:="1081";
                when 1082 => b:="1082";
                when 1083 => b:="1083";
                when 1084 => b:="1084";
                when 1085 => b:="1085";
                when 1086 => b:="1086";
                when 1087 => b:="1087";
                when 1088 => b:="1088";
                when 1089 => b:="1089";
                when 1090 => b:="1090";
                when 1091 => b:="1091";
                when 1092 => b:="1092";
                when 1093 => b:="1093";
                when 1094 => b:="1094";
                when 1095 => b:="1095";
                when 1096 => b:="1096";
                when 1097 => b:="1097";
                when 1098 => b:="1098";
                when 1099 => b:="1099";
                when 1100 => b:="1100";
                when 1101 => b:="1101";
                when 1102 => b:="1102";
                when 1103 => b:="1103";
                when 1104 => b:="1104";
                when 1105 => b:="1105";
                when 1106 => b:="1106";
                when 1107 => b:="1107";
                when 1108 => b:="1108";
                when 1109 => b:="1109";
                when 1110 => b:="1110";
                when 1111 => b:="1111";
                when 1112 => b:="1112";
                when 1113 => b:="1113";
                when 1114 => b:="1114";
                when 1115 => b:="1115";
                when 1116 => b:="1116";
                when 1117 => b:="1117";
                when 1118 => b:="1118";
                when 1119 => b:="1119";
                when 1120 => b:="1120";
                when 1121 => b:="1121";
                when 1122 => b:="1122";
                when 1123 => b:="1123";
                when 1124 => b:="1124";
                when 1125 => b:="1125";
                when 1126 => b:="1126";
                when 1127 => b:="1127";
                when 1128 => b:="1128";
                when 1129 => b:="1129";
                when 1130 => b:="1130";
                when 1131 => b:="1131";
                when 1132 => b:="1132";
                when 1133 => b:="1133";
                when 1134 => b:="1134";
                when 1135 => b:="1135";
                when 1136 => b:="1136";
                when 1137 => b:="1137";
                when 1138 => b:="1138";
                when 1139 => b:="1139";
                when 1140 => b:="1140";
                when 1141 => b:="1141";
                when 1142 => b:="1142";
                when 1143 => b:="1143";
                when 1144 => b:="1144";
                when 1145 => b:="1145";
                when 1146 => b:="1146";
                when 1147 => b:="1147";
                when 1148 => b:="1148";
                when 1149 => b:="1149";
                when 1150 => b:="1150";
                when 1151 => b:="1151";
                when 1152 => b:="1152";
                when 1153 => b:="1153";
                when 1154 => b:="1154";
                when 1155 => b:="1155";
                when 1156 => b:="1156";
                when 1157 => b:="1157";
                when 1158 => b:="1158";
                when 1159 => b:="1159";
                when 1160 => b:="1160";
                when 1161 => b:="1161";
                when 1162 => b:="1162";
                when 1163 => b:="1163";
                when 1164 => b:="1164";
                when 1165 => b:="1165";
                when 1166 => b:="1166";
                when 1167 => b:="1167";
                when 1168 => b:="1168";
                when 1169 => b:="1169";
                when 1170 => b:="1170";
                when 1171 => b:="1171";
                when 1172 => b:="1172";
                when 1173 => b:="1173";
                when 1174 => b:="1174";
                when 1175 => b:="1175";
                when 1176 => b:="1176";
                when 1177 => b:="1177";
                when 1178 => b:="1178";
                when 1179 => b:="1179";
                when 1180 => b:="1180";
                when 1181 => b:="1181";
                when 1182 => b:="1182";
                when 1183 => b:="1183";
                when 1184 => b:="1184";
                when 1185 => b:="1185";
                when 1186 => b:="1186";
                when 1187 => b:="1187";
                when 1188 => b:="1188";
                when 1189 => b:="1189";
                when 1190 => b:="1190";
                when 1191 => b:="1191";
                when 1192 => b:="1192";
                when 1193 => b:="1193";
                when 1194 => b:="1194";
                when 1195 => b:="1195";
                when 1196 => b:="1196";
                when 1197 => b:="1197";
                when 1198 => b:="1198";
                when 1199 => b:="1199";
                when 1200 => b:="1200";
                when 1201 => b:="1201";
                when 1202 => b:="1202";
                when 1203 => b:="1203";
                when 1204 => b:="1204";
                when 1205 => b:="1205";
                when 1206 => b:="1206";
                when 1207 => b:="1207";
                when 1208 => b:="1208";
                when 1209 => b:="1209";
                when 1210 => b:="1210";
                when 1211 => b:="1211";
                when 1212 => b:="1212";
                when 1213 => b:="1213";
                when 1214 => b:="1214";
                when 1215 => b:="1215";
                when 1216 => b:="1216";
                when 1217 => b:="1217";
                when 1218 => b:="1218";
                when 1219 => b:="1219";
                when 1220 => b:="1220";
                when 1221 => b:="1221";
                when 1222 => b:="1222";
                when 1223 => b:="1223";
                when 1224 => b:="1224";
                when 1225 => b:="1225";
                when 1226 => b:="1226";
                when 1227 => b:="1227";
                when 1228 => b:="1228";
                when 1229 => b:="1229";
                when 1230 => b:="1230";
                when 1231 => b:="1231";
                when 1232 => b:="1232";
                when 1233 => b:="1233";
                when 1234 => b:="1234";
                when 1235 => b:="1235";
                when 1236 => b:="1236";
                when 1237 => b:="1237";
                when 1238 => b:="1238";
                when 1239 => b:="1239";
                when 1240 => b:="1240";
                when 1241 => b:="1241";
                when 1242 => b:="1242";
                when 1243 => b:="1243";
                when 1244 => b:="1244";
                when 1245 => b:="1245";
                when 1246 => b:="1246";
                when 1247 => b:="1247";
                when 1248 => b:="1248";
                when 1249 => b:="1249";
                when 1250 => b:="1250";
                when 1251 => b:="1251";
                when 1252 => b:="1252";
                when 1253 => b:="1253";
                when 1254 => b:="1254";
                when 1255 => b:="1255";
                when 1256 => b:="1256";
                when 1257 => b:="1257";
                when 1258 => b:="1258";
                when 1259 => b:="1259";
                when 1260 => b:="1260";
                when 1261 => b:="1261";
                when 1262 => b:="1262";
                when 1263 => b:="1263";
                when 1264 => b:="1264";
                when 1265 => b:="1265";
                when 1266 => b:="1266";
                when 1267 => b:="1267";
                when 1268 => b:="1268";
                when 1269 => b:="1269";
                when 1270 => b:="1270";
                when 1271 => b:="1271";
                when 1272 => b:="1272";
                when 1273 => b:="1273";
                when 1274 => b:="1274";
                when 1275 => b:="1275";
                when 1276 => b:="1276";
                when 1277 => b:="1277";
                when 1278 => b:="1278";
                when 1279 => b:="1279";
                when 1280 => b:="1280";
                when 1281 => b:="1281";
                when 1282 => b:="1282";
                when 1283 => b:="1283";
                when 1284 => b:="1284";
                when 1285 => b:="1285";
                when 1286 => b:="1286";
                when 1287 => b:="1287";
                when 1288 => b:="1288";
                when 1289 => b:="1289";
                when 1290 => b:="1290";
                when 1291 => b:="1291";
                when 1292 => b:="1292";
                when 1293 => b:="1293";
                when 1294 => b:="1294";
                when 1295 => b:="1295";
                when 1296 => b:="1296";
                when 1297 => b:="1297";
                when 1298 => b:="1298";
                when 1299 => b:="1299";
                when 1300 => b:="1300";
                when 1301 => b:="1301";
                when 1302 => b:="1302";
                when 1303 => b:="1303";
                when 1304 => b:="1304";
                when 1305 => b:="1305";
                when 1306 => b:="1306";
                when 1307 => b:="1307";
                when 1308 => b:="1308";
                when 1309 => b:="1309";
                when 1310 => b:="1310";
                when 1311 => b:="1311";
                when 1312 => b:="1312";
                when 1313 => b:="1313";
                when 1314 => b:="1314";
                when 1315 => b:="1315";
                when 1316 => b:="1316";
                when 1317 => b:="1317";
                when 1318 => b:="1318";
                when 1319 => b:="1319";
                when 1320 => b:="1320";
                when 1321 => b:="1321";
                when 1322 => b:="1322";
                when 1323 => b:="1323";
                when 1324 => b:="1324";
                when 1325 => b:="1325";
                when 1326 => b:="1326";
                when 1327 => b:="1327";
                when 1328 => b:="1328";
                when 1329 => b:="1329";
                when 1330 => b:="1330";
                when 1331 => b:="1331";
                when 1332 => b:="1332";
                when 1333 => b:="1333";
                when 1334 => b:="1334";
                when 1335 => b:="1335";
                when 1336 => b:="1336";
                when 1337 => b:="1337";
                when 1338 => b:="1338";
                when 1339 => b:="1339";
                when 1340 => b:="1340";
                when 1341 => b:="1341";
                when 1342 => b:="1342";
                when 1343 => b:="1343";
                when 1344 => b:="1344";
                when 1345 => b:="1345";
                when 1346 => b:="1346";
                when 1347 => b:="1347";
                when 1348 => b:="1348";
                when 1349 => b:="1349";
                when 1350 => b:="1350";
                when 1351 => b:="1351";
                when 1352 => b:="1352";
                when 1353 => b:="1353";
                when 1354 => b:="1354";
                when 1355 => b:="1355";
                when 1356 => b:="1356";
                when 1357 => b:="1357";
                when 1358 => b:="1358";
                when 1359 => b:="1359";
                when 1360 => b:="1360";
                when 1361 => b:="1361";
                when 1362 => b:="1362";
                when 1363 => b:="1363";
                when 1364 => b:="1364";
                when 1365 => b:="1365";
                when 1366 => b:="1366";
                when 1367 => b:="1367";
                when 1368 => b:="1368";
                when 1369 => b:="1369";
                when 1370 => b:="1370";
                when 1371 => b:="1371";
                when 1372 => b:="1372";
                when 1373 => b:="1373";
                when 1374 => b:="1374";
                when 1375 => b:="1375";
                when 1376 => b:="1376";
                when 1377 => b:="1377";
                when 1378 => b:="1378";
                when 1379 => b:="1379";
                when 1380 => b:="1380";
                when 1381 => b:="1381";
                when 1382 => b:="1382";
                when 1383 => b:="1383";
                when 1384 => b:="1384";
                when 1385 => b:="1385";
                when 1386 => b:="1386";
                when 1387 => b:="1387";
                when 1388 => b:="1388";
                when 1389 => b:="1389";
                when 1390 => b:="1390";
                when 1391 => b:="1391";
                when 1392 => b:="1392";
                when 1393 => b:="1393";
                when 1394 => b:="1394";
                when 1395 => b:="1395";
                when 1396 => b:="1396";
                when 1397 => b:="1397";
                when 1398 => b:="1398";
                when 1399 => b:="1399";
                when 1400 => b:="1400";
                when 1401 => b:="1401";
                when 1402 => b:="1402";
                when 1403 => b:="1403";
                when 1404 => b:="1404";
                when 1405 => b:="1405";
                when 1406 => b:="1406";
                when 1407 => b:="1407";
                when 1408 => b:="1408";
                when 1409 => b:="1409";
                when 1410 => b:="1410";
                when 1411 => b:="1411";
                when 1412 => b:="1412";
                when 1413 => b:="1413";
                when 1414 => b:="1414";
                when 1415 => b:="1415";
                when 1416 => b:="1416";
                when 1417 => b:="1417";
                when 1418 => b:="1418";
                when 1419 => b:="1419";
                when 1420 => b:="1420";
                when 1421 => b:="1421";
                when 1422 => b:="1422";
                when 1423 => b:="1423";
                when 1424 => b:="1424";
                when 1425 => b:="1425";
                when 1426 => b:="1426";
                when 1427 => b:="1427";
                when 1428 => b:="1428";
                when 1429 => b:="1429";
                when 1430 => b:="1430";
                when 1431 => b:="1431";
                when 1432 => b:="1432";
                when 1433 => b:="1433";
                when 1434 => b:="1434";
                when 1435 => b:="1435";
                when 1436 => b:="1436";
                when 1437 => b:="1437";
                when 1438 => b:="1438";
                when 1439 => b:="1439";
                when 1440 => b:="1440";
                when 1441 => b:="1441";
                when 1442 => b:="1442";
                when 1443 => b:="1443";
                when 1444 => b:="1444";
                when 1445 => b:="1445";
                when 1446 => b:="1446";
                when 1447 => b:="1447";
                when 1448 => b:="1448";
                when 1449 => b:="1449";
                when 1450 => b:="1450";
                when 1451 => b:="1451";
                when 1452 => b:="1452";
                when 1453 => b:="1453";
                when 1454 => b:="1454";
                when 1455 => b:="1455";
                when 1456 => b:="1456";
                when 1457 => b:="1457";
                when 1458 => b:="1458";
                when 1459 => b:="1459";
                when 1460 => b:="1460";
                when 1461 => b:="1461";
                when 1462 => b:="1462";
                when 1463 => b:="1463";
                when 1464 => b:="1464";
                when 1465 => b:="1465";
                when 1466 => b:="1466";
                when 1467 => b:="1467";
                when 1468 => b:="1468";
                when 1469 => b:="1469";
                when 1470 => b:="1470";
                when 1471 => b:="1471";
                when 1472 => b:="1472";
                when 1473 => b:="1473";
                when 1474 => b:="1474";
                when 1475 => b:="1475";
                when 1476 => b:="1476";
                when 1477 => b:="1477";
                when 1478 => b:="1478";
                when 1479 => b:="1479";
                when 1480 => b:="1480";
                when 1481 => b:="1481";
                when 1482 => b:="1482";
                when 1483 => b:="1483";
                when 1484 => b:="1484";
                when 1485 => b:="1485";
                when 1486 => b:="1486";
                when 1487 => b:="1487";
                when 1488 => b:="1488";
                when 1489 => b:="1489";
                when 1490 => b:="1490";
                when 1491 => b:="1491";
                when 1492 => b:="1492";
                when 1493 => b:="1493";
                when 1494 => b:="1494";
                when 1495 => b:="1495";
                when 1496 => b:="1496";
                when 1497 => b:="1497";
                when 1498 => b:="1498";
                when 1499 => b:="1499";
                when 1500 => b:="1500";
                when 1501 => b:="1501";
                when 1502 => b:="1502";
                when 1503 => b:="1503";
                when 1504 => b:="1504";
                when 1505 => b:="1505";
                when 1506 => b:="1506";
                when 1507 => b:="1507";
                when 1508 => b:="1508";
                when 1509 => b:="1509";
                when 1510 => b:="1510";
                when 1511 => b:="1511";
                when 1512 => b:="1512";
                when 1513 => b:="1513";
                when 1514 => b:="1514";
                when 1515 => b:="1515";
                when 1516 => b:="1516";
                when 1517 => b:="1517";
                when 1518 => b:="1518";
                when 1519 => b:="1519";
                when 1520 => b:="1520";
                when 1521 => b:="1521";
                when 1522 => b:="1522";
                when 1523 => b:="1523";
                when 1524 => b:="1524";
                when 1525 => b:="1525";
                when 1526 => b:="1526";
                when 1527 => b:="1527";
                when 1528 => b:="1528";
                when 1529 => b:="1529";
                when 1530 => b:="1530";
                when 1531 => b:="1531";
                when 1532 => b:="1532";
                when 1533 => b:="1533";
                when 1534 => b:="1534";
                when 1535 => b:="1535";
                when 1536 => b:="1536";
                when 1537 => b:="1537";
                when 1538 => b:="1538";
                when 1539 => b:="1539";
                when 1540 => b:="1540";
                when 1541 => b:="1541";
                when 1542 => b:="1542";
                when 1543 => b:="1543";
                when 1544 => b:="1544";
                when 1545 => b:="1545";
                when 1546 => b:="1546";
                when 1547 => b:="1547";
                when 1548 => b:="1548";
                when 1549 => b:="1549";
                when 1550 => b:="1550";
                when 1551 => b:="1551";
                when 1552 => b:="1552";
                when 1553 => b:="1553";
                when 1554 => b:="1554";
                when 1555 => b:="1555";
                when 1556 => b:="1556";
                when 1557 => b:="1557";
                when 1558 => b:="1558";
                when 1559 => b:="1559";
                when 1560 => b:="1560";
                when 1561 => b:="1561";
                when 1562 => b:="1562";
                when 1563 => b:="1563";
                when 1564 => b:="1564";
                when 1565 => b:="1565";
                when 1566 => b:="1566";
                when 1567 => b:="1567";
                when 1568 => b:="1568";
                when 1569 => b:="1569";
                when 1570 => b:="1570";
                when 1571 => b:="1571";
                when 1572 => b:="1572";
                when 1573 => b:="1573";
                when 1574 => b:="1574";
                when 1575 => b:="1575";
                when 1576 => b:="1576";
                when 1577 => b:="1577";
                when 1578 => b:="1578";
                when 1579 => b:="1579";
                when 1580 => b:="1580";
                when 1581 => b:="1581";
                when 1582 => b:="1582";
                when 1583 => b:="1583";
                when 1584 => b:="1584";
                when 1585 => b:="1585";
                when 1586 => b:="1586";
                when 1587 => b:="1587";
                when 1588 => b:="1588";
                when 1589 => b:="1589";
                when 1590 => b:="1590";
                when 1591 => b:="1591";
                when 1592 => b:="1592";
                when 1593 => b:="1593";
                when 1594 => b:="1594";
                when 1595 => b:="1595";
                when 1596 => b:="1596";
                when 1597 => b:="1597";
                when 1598 => b:="1598";
                when 1599 => b:="1599";
                when 1600 => b:="1600";
                when 1601 => b:="1601";
                when 1602 => b:="1602";
                when 1603 => b:="1603";
                when 1604 => b:="1604";
                when 1605 => b:="1605";
                when 1606 => b:="1606";
                when 1607 => b:="1607";
                when 1608 => b:="1608";
                when 1609 => b:="1609";
                when 1610 => b:="1610";
                when 1611 => b:="1611";
                when 1612 => b:="1612";
                when 1613 => b:="1613";
                when 1614 => b:="1614";
                when 1615 => b:="1615";
                when 1616 => b:="1616";
                when 1617 => b:="1617";
                when 1618 => b:="1618";
                when 1619 => b:="1619";
                when 1620 => b:="1620";
                when 1621 => b:="1621";
                when 1622 => b:="1622";
                when 1623 => b:="1623";
                when 1624 => b:="1624";
                when 1625 => b:="1625";
                when 1626 => b:="1626";
                when 1627 => b:="1627";
                when 1628 => b:="1628";
                when 1629 => b:="1629";
                when 1630 => b:="1630";
                when 1631 => b:="1631";
                when 1632 => b:="1632";
                when 1633 => b:="1633";
                when 1634 => b:="1634";
                when 1635 => b:="1635";
                when 1636 => b:="1636";
                when 1637 => b:="1637";
                when 1638 => b:="1638";
                when 1639 => b:="1639";
                when 1640 => b:="1640";
                when 1641 => b:="1641";
                when 1642 => b:="1642";
                when 1643 => b:="1643";
                when 1644 => b:="1644";
                when 1645 => b:="1645";
                when 1646 => b:="1646";
                when 1647 => b:="1647";
                when 1648 => b:="1648";
                when 1649 => b:="1649";
                when 1650 => b:="1650";
                when 1651 => b:="1651";
                when 1652 => b:="1652";
                when 1653 => b:="1653";
                when 1654 => b:="1654";
                when 1655 => b:="1655";
                when 1656 => b:="1656";
                when 1657 => b:="1657";
                when 1658 => b:="1658";
                when 1659 => b:="1659";
                when 1660 => b:="1660";
                when 1661 => b:="1661";
                when 1662 => b:="1662";
                when 1663 => b:="1663";
                when 1664 => b:="1664";
                when 1665 => b:="1665";
                when 1666 => b:="1666";
                when 1667 => b:="1667";
                when 1668 => b:="1668";
                when 1669 => b:="1669";
                when 1670 => b:="1670";
                when 1671 => b:="1671";
                when 1672 => b:="1672";
                when 1673 => b:="1673";
                when 1674 => b:="1674";
                when 1675 => b:="1675";
                when 1676 => b:="1676";
                when 1677 => b:="1677";
                when 1678 => b:="1678";
                when 1679 => b:="1679";
                when 1680 => b:="1680";
                when 1681 => b:="1681";
                when 1682 => b:="1682";
                when 1683 => b:="1683";
                when 1684 => b:="1684";
                when 1685 => b:="1685";
                when 1686 => b:="1686";
                when 1687 => b:="1687";
                when 1688 => b:="1688";
                when 1689 => b:="1689";
                when 1690 => b:="1690";
                when 1691 => b:="1691";
                when 1692 => b:="1692";
                when 1693 => b:="1693";
                when 1694 => b:="1694";
                when 1695 => b:="1695";
                when 1696 => b:="1696";
                when 1697 => b:="1697";
                when 1698 => b:="1698";
                when 1699 => b:="1699";
                when 1700 => b:="1700";
                when 1701 => b:="1701";
                when 1702 => b:="1702";
                when 1703 => b:="1703";
                when 1704 => b:="1704";
                when 1705 => b:="1705";
                when 1706 => b:="1706";
                when 1707 => b:="1707";
                when 1708 => b:="1708";
                when 1709 => b:="1709";
                when 1710 => b:="1710";
                when 1711 => b:="1711";
                when 1712 => b:="1712";
                when 1713 => b:="1713";
                when 1714 => b:="1714";
                when 1715 => b:="1715";
                when 1716 => b:="1716";
                when 1717 => b:="1717";
                when 1718 => b:="1718";
                when 1719 => b:="1719";
                when 1720 => b:="1720";
                when 1721 => b:="1721";
                when 1722 => b:="1722";
                when 1723 => b:="1723";
                when 1724 => b:="1724";
                when 1725 => b:="1725";
                when 1726 => b:="1726";
                when 1727 => b:="1727";
                when 1728 => b:="1728";
                when 1729 => b:="1729";
                when 1730 => b:="1730";
                when 1731 => b:="1731";
                when 1732 => b:="1732";
                when 1733 => b:="1733";
                when 1734 => b:="1734";
                when 1735 => b:="1735";
                when 1736 => b:="1736";
                when 1737 => b:="1737";
                when 1738 => b:="1738";
                when 1739 => b:="1739";
                when 1740 => b:="1740";
                when 1741 => b:="1741";
                when 1742 => b:="1742";
                when 1743 => b:="1743";
                when 1744 => b:="1744";
                when 1745 => b:="1745";
                when 1746 => b:="1746";
                when 1747 => b:="1747";
                when 1748 => b:="1748";
                when 1749 => b:="1749";
                when 1750 => b:="1750";
                when 1751 => b:="1751";
                when 1752 => b:="1752";
                when 1753 => b:="1753";
                when 1754 => b:="1754";
                when 1755 => b:="1755";
                when 1756 => b:="1756";
                when 1757 => b:="1757";
                when 1758 => b:="1758";
                when 1759 => b:="1759";
                when 1760 => b:="1760";
                when 1761 => b:="1761";
                when 1762 => b:="1762";
                when 1763 => b:="1763";
                when 1764 => b:="1764";
                when 1765 => b:="1765";
                when 1766 => b:="1766";
                when 1767 => b:="1767";
                when 1768 => b:="1768";
                when 1769 => b:="1769";
                when 1770 => b:="1770";
                when 1771 => b:="1771";
                when 1772 => b:="1772";
                when 1773 => b:="1773";
                when 1774 => b:="1774";
                when 1775 => b:="1775";
                when 1776 => b:="1776";
                when 1777 => b:="1777";
                when 1778 => b:="1778";
                when 1779 => b:="1779";
                when 1780 => b:="1780";
                when 1781 => b:="1781";
                when 1782 => b:="1782";
                when 1783 => b:="1783";
                when 1784 => b:="1784";
                when 1785 => b:="1785";
                when 1786 => b:="1786";
                when 1787 => b:="1787";
                when 1788 => b:="1788";
                when 1789 => b:="1789";
                when 1790 => b:="1790";
                when 1791 => b:="1791";
                when 1792 => b:="1792";
                when 1793 => b:="1793";
                when 1794 => b:="1794";
                when 1795 => b:="1795";
                when 1796 => b:="1796";
                when 1797 => b:="1797";
                when 1798 => b:="1798";
                when 1799 => b:="1799";
                when 1800 => b:="1800";
                when 1801 => b:="1801";
                when 1802 => b:="1802";
                when 1803 => b:="1803";
                when 1804 => b:="1804";
                when 1805 => b:="1805";
                when 1806 => b:="1806";
                when 1807 => b:="1807";
                when 1808 => b:="1808";
                when 1809 => b:="1809";
                when 1810 => b:="1810";
                when 1811 => b:="1811";
                when 1812 => b:="1812";
                when 1813 => b:="1813";
                when 1814 => b:="1814";
                when 1815 => b:="1815";
                when 1816 => b:="1816";
                when 1817 => b:="1817";
                when 1818 => b:="1818";
                when 1819 => b:="1819";
                when 1820 => b:="1820";
                when 1821 => b:="1821";
                when 1822 => b:="1822";
                when 1823 => b:="1823";
                when 1824 => b:="1824";
                when 1825 => b:="1825";
                when 1826 => b:="1826";
                when 1827 => b:="1827";
                when 1828 => b:="1828";
                when 1829 => b:="1829";
                when 1830 => b:="1830";
                when 1831 => b:="1831";
                when 1832 => b:="1832";
                when 1833 => b:="1833";
                when 1834 => b:="1834";
                when 1835 => b:="1835";
                when 1836 => b:="1836";
                when 1837 => b:="1837";
                when 1838 => b:="1838";
                when 1839 => b:="1839";
                when 1840 => b:="1840";
                when 1841 => b:="1841";
                when 1842 => b:="1842";
                when 1843 => b:="1843";
                when 1844 => b:="1844";
                when 1845 => b:="1845";
                when 1846 => b:="1846";
                when 1847 => b:="1847";
                when 1848 => b:="1848";
                when 1849 => b:="1849";
                when 1850 => b:="1850";
                when 1851 => b:="1851";
                when 1852 => b:="1852";
                when 1853 => b:="1853";
                when 1854 => b:="1854";
                when 1855 => b:="1855";
                when 1856 => b:="1856";
                when 1857 => b:="1857";
                when 1858 => b:="1858";
                when 1859 => b:="1859";
                when 1860 => b:="1860";
                when 1861 => b:="1861";
                when 1862 => b:="1862";
                when 1863 => b:="1863";
                when 1864 => b:="1864";
                when 1865 => b:="1865";
                when 1866 => b:="1866";
                when 1867 => b:="1867";
                when 1868 => b:="1868";
                when 1869 => b:="1869";
                when 1870 => b:="1870";
                when 1871 => b:="1871";
                when 1872 => b:="1872";
                when 1873 => b:="1873";
                when 1874 => b:="1874";
                when 1875 => b:="1875";
                when 1876 => b:="1876";
                when 1877 => b:="1877";
                when 1878 => b:="1878";
                when 1879 => b:="1879";
                when 1880 => b:="1880";
                when 1881 => b:="1881";
                when 1882 => b:="1882";
                when 1883 => b:="1883";
                when 1884 => b:="1884";
                when 1885 => b:="1885";
                when 1886 => b:="1886";
                when 1887 => b:="1887";
                when 1888 => b:="1888";
                when 1889 => b:="1889";
                when 1890 => b:="1890";
                when 1891 => b:="1891";
                when 1892 => b:="1892";
                when 1893 => b:="1893";
                when 1894 => b:="1894";
                when 1895 => b:="1895";
                when 1896 => b:="1896";
                when 1897 => b:="1897";
                when 1898 => b:="1898";
                when 1899 => b:="1899";
                when 1900 => b:="1900";
                when 1901 => b:="1901";
                when 1902 => b:="1902";
                when 1903 => b:="1903";
                when 1904 => b:="1904";
                when 1905 => b:="1905";
                when 1906 => b:="1906";
                when 1907 => b:="1907";
                when 1908 => b:="1908";
                when 1909 => b:="1909";
                when 1910 => b:="1910";
                when 1911 => b:="1911";
                when 1912 => b:="1912";
                when 1913 => b:="1913";
                when 1914 => b:="1914";
                when 1915 => b:="1915";
                when 1916 => b:="1916";
                when 1917 => b:="1917";
                when 1918 => b:="1918";
                when 1919 => b:="1919";
                when 1920 => b:="1920";
                when 1921 => b:="1921";
                when 1922 => b:="1922";
                when 1923 => b:="1923";
                when 1924 => b:="1924";
                when 1925 => b:="1925";
                when 1926 => b:="1926";
                when 1927 => b:="1927";
                when 1928 => b:="1928";
                when 1929 => b:="1929";
                when 1930 => b:="1930";
                when 1931 => b:="1931";
                when 1932 => b:="1932";
                when 1933 => b:="1933";
                when 1934 => b:="1934";
                when 1935 => b:="1935";
                when 1936 => b:="1936";
                when 1937 => b:="1937";
                when 1938 => b:="1938";
                when 1939 => b:="1939";
                when 1940 => b:="1940";
                when 1941 => b:="1941";
                when 1942 => b:="1942";
                when 1943 => b:="1943";
                when 1944 => b:="1944";
                when 1945 => b:="1945";
                when 1946 => b:="1946";
                when 1947 => b:="1947";
                when 1948 => b:="1948";
                when 1949 => b:="1949";
                when 1950 => b:="1950";
                when 1951 => b:="1951";
                when 1952 => b:="1952";
                when 1953 => b:="1953";
                when 1954 => b:="1954";
                when 1955 => b:="1955";
                when 1956 => b:="1956";
                when 1957 => b:="1957";
                when 1958 => b:="1958";
                when 1959 => b:="1959";
                when 1960 => b:="1960";
                when 1961 => b:="1961";
                when 1962 => b:="1962";
                when 1963 => b:="1963";
                when 1964 => b:="1964";
                when 1965 => b:="1965";
                when 1966 => b:="1966";
                when 1967 => b:="1967";
                when 1968 => b:="1968";
                when 1969 => b:="1969";
                when 1970 => b:="1970";
                when 1971 => b:="1971";
                when 1972 => b:="1972";
                when 1973 => b:="1973";
                when 1974 => b:="1974";
                when 1975 => b:="1975";
                when 1976 => b:="1976";
                when 1977 => b:="1977";
                when 1978 => b:="1978";
                when 1979 => b:="1979";
                when 1980 => b:="1980";
                when 1981 => b:="1981";
                when 1982 => b:="1982";
                when 1983 => b:="1983";
                when 1984 => b:="1984";
                when 1985 => b:="1985";
                when 1986 => b:="1986";
                when 1987 => b:="1987";
                when 1988 => b:="1988";
                when 1989 => b:="1989";
                when 1990 => b:="1990";
                when 1991 => b:="1991";
                when 1992 => b:="1992";
                when 1993 => b:="1993";
                when 1994 => b:="1994";
                when 1995 => b:="1995";
                when 1996 => b:="1996";
                when 1997 => b:="1997";
                when 1998 => b:="1998";
                when 2000 => b:="2000";
                when 2001 => b:="2001";
                when 2002 => b:="2002";
                when 2003 => b:="2003";
                when 2004 => b:="2004";
                when 2005 => b:="2005";
                when 2006 => b:="2006";
                when 2007 => b:="2007";
                when 2008 => b:="2008";
                when 2009 => b:="2009";
                when 2010 => b:="2010";
                when 2011 => b:="2011";
                when 2012 => b:="2012";
                when 2013 => b:="2013";
                when 2014 => b:="2014";
                when 2015 => b:="2015";
                when 2016 => b:="2016";
                when 2017 => b:="2017";
                when 2018 => b:="2018";
                when 2019 => b:="2019";
                when 2020 => b:="2020";
                when 2021 => b:="2021";
                when 2022 => b:="2022";
                when 2023 => b:="2023";
                when 2024 => b:="2024";
                when 2025 => b:="2025";
                when 2026 => b:="2026";
                when 2027 => b:="2027";
                when 2028 => b:="2028";
                when 2029 => b:="2029";
                when 2030 => b:="2030";
                when 2031 => b:="2031";
                when 2032 => b:="2032";
                when 2033 => b:="2033";
                when 2034 => b:="2034";
                when 2035 => b:="2035";
                when 2036 => b:="2036";
                when 2037 => b:="2037";
                when 2038 => b:="2038";
                when 2039 => b:="2039";
                when 2040 => b:="2040";
                when 2041 => b:="2041";
                when 2042 => b:="2042";
                when 2043 => b:="2043";
                when 2044 => b:="2044";
                when 2045 => b:="2045";
                when 2046 => b:="2046";
                when 2047 => b:="2047";
                when 2048 => b:="2048";
                when 2049 => b:="2049";
                when 2050 => b:="2050";
                when 2051 => b:="2051";
                when 2052 => b:="2052";
                when 2053 => b:="2053";
                when 2054 => b:="2054";
                when 2055 => b:="2055";
                when 2056 => b:="2056";
                when 2057 => b:="2057";
                when 2058 => b:="2058";
                when 2059 => b:="2059";
                when 2060 => b:="2060";
                when 2061 => b:="2061";
                when 2062 => b:="2062";
                when 2063 => b:="2063";
                when 2064 => b:="2064";
                when 2065 => b:="2065";
                when 2066 => b:="2066";
                when 2067 => b:="2067";
                when 2068 => b:="2068";
                when 2069 => b:="2069";
                when 2070 => b:="2070";
                when 2071 => b:="2071";
                when 2072 => b:="2072";
                when 2073 => b:="2073";
                when 2074 => b:="2074";
                when 2075 => b:="2075";
                when 2076 => b:="2076";
                when 2077 => b:="2077";
                when 2078 => b:="2078";
                when 2079 => b:="2079";
                when 2080 => b:="2080";
                when 2081 => b:="2081";
                when 2082 => b:="2082";
                when 2083 => b:="2083";
                when 2084 => b:="2084";
                when 2085 => b:="2085";
                when 2086 => b:="2086";
                when 2087 => b:="2087";
                when 2088 => b:="2088";
                when 2089 => b:="2089";
                when 2090 => b:="2090";
                when 2091 => b:="2091";
                when 2092 => b:="2092";
                when 2093 => b:="2093";
                when 2094 => b:="2094";
                when 2095 => b:="2095";
                when 2096 => b:="2096";
                when 2097 => b:="2097";
                when 2098 => b:="2098";
                when 2099 => b:="2099";
                when 2100 => b:="2100";
                when 2101 => b:="2101";
                when 2102 => b:="2102";
                when 2103 => b:="2103";
                when 2104 => b:="2104";
                when 2105 => b:="2105";
                when 2106 => b:="2106";
                when 2107 => b:="2107";
                when 2108 => b:="2108";
                when 2109 => b:="2109";
                when 2110 => b:="2110";
                when 2111 => b:="2111";
                when 2112 => b:="2112";
                when 2113 => b:="2113";
                when 2114 => b:="2114";
                when 2115 => b:="2115";
                when 2116 => b:="2116";
                when 2117 => b:="2117";
                when 2118 => b:="2118";
                when 2119 => b:="2119";
                when 2120 => b:="2120";
                when 2121 => b:="2121";
                when 2122 => b:="2122";
                when 2123 => b:="2123";
                when 2124 => b:="2124";
                when 2125 => b:="2125";
                when 2126 => b:="2126";
                when 2127 => b:="2127";
                when 2128 => b:="2128";
                when 2129 => b:="2129";
                when 2130 => b:="2130";
                when 2131 => b:="2131";
                when 2132 => b:="2132";
                when 2133 => b:="2133";
                when 2134 => b:="2134";
                when 2135 => b:="2135";
                when 2136 => b:="2136";
                when 2137 => b:="2137";
                when 2138 => b:="2138";
                when 2139 => b:="2139";
                when 2140 => b:="2140";
                when 2141 => b:="2141";
                when 2142 => b:="2142";
                when 2143 => b:="2143";
                when 2144 => b:="2144";
                when 2145 => b:="2145";
                when 2146 => b:="2146";
                when 2147 => b:="2147";
                when 2148 => b:="2148";
                when 2149 => b:="2149";
                when 2150 => b:="2150";
                when 2151 => b:="2151";
                when 2152 => b:="2152";
                when 2153 => b:="2153";
                when 2154 => b:="2154";
                when 2155 => b:="2155";
                when 2156 => b:="2156";
                when 2157 => b:="2157";
                when 2158 => b:="2158";
                when 2159 => b:="2159";
                when 2160 => b:="2160";
                when 2161 => b:="2161";
                when 2162 => b:="2162";
                when 2163 => b:="2163";
                when 2164 => b:="2164";
                when 2165 => b:="2165";
                when 2166 => b:="2166";
                when 2167 => b:="2167";
                when 2168 => b:="2168";
                when 2169 => b:="2169";
                when 2170 => b:="2170";
                when 2171 => b:="2171";
                when 2172 => b:="2172";
                when 2173 => b:="2173";
                when 2174 => b:="2174";
                when 2175 => b:="2175";
                when 2176 => b:="2176";
                when 2177 => b:="2177";
                when 2178 => b:="2178";
                when 2179 => b:="2179";
                when 2180 => b:="2180";
                when 2181 => b:="2181";
                when 2182 => b:="2182";
                when 2183 => b:="2183";
                when 2184 => b:="2184";
                when 2185 => b:="2185";
                when 2186 => b:="2186";
                when 2187 => b:="2187";
                when 2188 => b:="2188";
                when 2189 => b:="2189";
                when 2190 => b:="2190";
                when 2191 => b:="2191";
                when 2192 => b:="2192";
                when 2193 => b:="2193";
                when 2194 => b:="2194";
                when 2195 => b:="2195";
                when 2196 => b:="2196";
                when 2197 => b:="2197";
                when 2198 => b:="2198";
                when 2199 => b:="2199";
                when 2200 => b:="2200";
                when 2201 => b:="2201";
                when 2202 => b:="2202";
                when 2203 => b:="2203";
                when 2204 => b:="2204";
                when 2205 => b:="2205";
                when 2206 => b:="2206";
                when 2207 => b:="2207";
                when 2208 => b:="2208";
                when 2209 => b:="2209";
                when 2210 => b:="2210";
                when 2211 => b:="2211";
                when 2212 => b:="2212";
                when 2213 => b:="2213";
                when 2214 => b:="2214";
                when 2215 => b:="2215";
                when 2216 => b:="2216";
                when 2217 => b:="2217";
                when 2218 => b:="2218";
                when 2219 => b:="2219";
                when 2220 => b:="2220";
                when 2221 => b:="2221";
                when 2222 => b:="2222";
                when 2223 => b:="2223";
                when 2224 => b:="2224";
                when 2225 => b:="2225";
                when 2226 => b:="2226";
                when 2227 => b:="2227";
                when 2228 => b:="2228";
                when 2229 => b:="2229";
                when 2230 => b:="2230";
                when 2231 => b:="2231";
                when 2232 => b:="2232";
                when 2233 => b:="2233";
                when 2234 => b:="2234";
                when 2235 => b:="2235";
                when 2236 => b:="2236";
                when 2237 => b:="2237";
                when 2238 => b:="2238";
                when 2239 => b:="2239";
                when 2240 => b:="2240";
                when 2241 => b:="2241";
                when 2242 => b:="2242";
                when 2243 => b:="2243";
                when 2244 => b:="2244";
                when 2245 => b:="2245";
                when 2246 => b:="2246";
                when 2247 => b:="2247";
                when 2248 => b:="2248";
                when 2249 => b:="2249";
                when 2250 => b:="2250";
                when 2251 => b:="2251";
                when 2252 => b:="2252";
                when 2253 => b:="2253";
                when 2254 => b:="2254";
                when 2255 => b:="2255";
                when 2256 => b:="2256";
                when 2257 => b:="2257";
                when 2258 => b:="2258";
                when 2259 => b:="2259";
                when 2260 => b:="2260";
                when 2261 => b:="2261";
                when 2262 => b:="2262";
                when 2263 => b:="2263";
                when 2264 => b:="2264";
                when 2265 => b:="2265";
                when 2266 => b:="2266";
                when 2267 => b:="2267";
                when 2268 => b:="2268";
                when 2269 => b:="2269";
                when 2270 => b:="2270";
                when 2271 => b:="2271";
                when 2272 => b:="2272";
                when 2273 => b:="2273";
                when 2274 => b:="2274";
                when 2275 => b:="2275";
                when 2276 => b:="2276";
                when 2277 => b:="2277";
                when 2278 => b:="2278";
                when 2279 => b:="2279";
                when 2280 => b:="2280";
                when 2281 => b:="2281";
                when 2282 => b:="2282";
                when 2283 => b:="2283";
                when 2284 => b:="2284";
                when 2285 => b:="2285";
                when 2286 => b:="2286";
                when 2287 => b:="2287";
                when 2288 => b:="2288";
                when 2289 => b:="2289";
                when 2290 => b:="2290";
                when 2291 => b:="2291";
                when 2292 => b:="2292";
                when 2293 => b:="2293";
                when 2294 => b:="2294";
                when 2295 => b:="2295";
                when 2296 => b:="2296";
                when 2297 => b:="2297";
                when 2298 => b:="2298";
                when 2299 => b:="2299";
                when 2300 => b:="2300";
                when 2301 => b:="2301";
                when 2302 => b:="2302";
                when 2303 => b:="2303";
                when 2304 => b:="2304";
                when 2305 => b:="2305";
                when 2306 => b:="2306";
                when 2307 => b:="2307";
                when 2308 => b:="2308";
                when 2309 => b:="2309";
                when 2310 => b:="2310";
                when 2311 => b:="2311";
                when 2312 => b:="2312";
                when 2313 => b:="2313";
                when 2314 => b:="2314";
                when 2315 => b:="2315";
                when 2316 => b:="2316";
                when 2317 => b:="2317";
                when 2318 => b:="2318";
                when 2319 => b:="2319";
                when 2320 => b:="2320";
                when 2321 => b:="2321";
                when 2322 => b:="2322";
                when 2323 => b:="2323";
                when 2324 => b:="2324";
                when 2325 => b:="2325";
                when 2326 => b:="2326";
                when 2327 => b:="2327";
                when 2328 => b:="2328";
                when 2329 => b:="2329";
                when 2330 => b:="2330";
                when 2331 => b:="2331";
                when 2332 => b:="2332";
                when 2333 => b:="2333";
                when 2334 => b:="2334";
                when 2335 => b:="2335";
                when 2336 => b:="2336";
                when 2337 => b:="2337";
                when 2338 => b:="2338";
                when 2339 => b:="2339";
                when 2340 => b:="2340";
                when 2341 => b:="2341";
                when 2342 => b:="2342";
                when 2343 => b:="2343";
                when 2344 => b:="2344";
                when 2345 => b:="2345";
                when 2346 => b:="2346";
                when 2347 => b:="2347";
                when 2348 => b:="2348";
                when 2349 => b:="2349";
                when 2350 => b:="2350";
                when 2351 => b:="2351";
                when 2352 => b:="2352";
                when 2353 => b:="2353";
                when 2354 => b:="2354";
                when 2355 => b:="2355";
                when 2356 => b:="2356";
                when 2357 => b:="2357";
                when 2358 => b:="2358";
                when 2359 => b:="2359";
                when 2360 => b:="2360";
                when 2361 => b:="2361";
                when 2362 => b:="2362";
                when 2363 => b:="2363";
                when 2364 => b:="2364";
                when 2365 => b:="2365";
                when 2366 => b:="2366";
                when 2367 => b:="2367";
                when 2368 => b:="2368";
                when 2369 => b:="2369";
                when 2370 => b:="2370";
                when 2371 => b:="2371";
                when 2372 => b:="2372";
                when 2373 => b:="2373";
                when 2374 => b:="2374";
                when 2375 => b:="2375";
                when 2376 => b:="2376";
                when 2377 => b:="2377";
                when 2378 => b:="2378";
                when 2379 => b:="2379";
                when 2380 => b:="2380";
                when 2381 => b:="2381";
                when 2382 => b:="2382";
                when 2383 => b:="2383";
                when 2384 => b:="2384";
                when 2385 => b:="2385";
                when 2386 => b:="2386";
                when 2387 => b:="2387";
                when 2388 => b:="2388";
                when 2389 => b:="2389";
                when 2390 => b:="2390";
                when 2391 => b:="2391";
                when 2392 => b:="2392";
                when 2393 => b:="2393";
                when 2394 => b:="2394";
                when 2395 => b:="2395";
                when 2396 => b:="2396";
                when 2397 => b:="2397";
                when 2398 => b:="2398";
                when 2399 => b:="2399";
                when 2400 => b:="2400";
                when 2401 => b:="2401";
                when 2402 => b:="2402";
                when 2403 => b:="2403";
                when 2404 => b:="2404";
                when 2405 => b:="2405";
                when 2406 => b:="2406";
                when 2407 => b:="2407";
                when 2408 => b:="2408";
                when 2409 => b:="2409";
                when 2410 => b:="2410";
                when 2411 => b:="2411";
                when 2412 => b:="2412";
                when 2413 => b:="2413";
                when 2414 => b:="2414";
                when 2415 => b:="2415";
                when 2416 => b:="2416";
                when 2417 => b:="2417";
                when 2418 => b:="2418";
                when 2419 => b:="2419";
                when 2420 => b:="2420";
                when 2421 => b:="2421";
                when 2422 => b:="2422";
                when 2423 => b:="2423";
                when 2424 => b:="2424";
                when 2425 => b:="2425";
                when 2426 => b:="2426";
                when 2427 => b:="2427";
                when 2428 => b:="2428";
                when 2429 => b:="2429";
                when 2430 => b:="2430";
                when 2431 => b:="2431";
                when 2432 => b:="2432";
                when 2433 => b:="2433";
                when 2434 => b:="2434";
                when 2435 => b:="2435";
                when 2436 => b:="2436";
                when 2437 => b:="2437";
                when 2438 => b:="2438";
                when 2439 => b:="2439";
                when 2440 => b:="2440";
                when 2441 => b:="2441";
                when 2442 => b:="2442";
                when 2443 => b:="2443";
                when 2444 => b:="2444";
                when 2445 => b:="2445";
                when 2446 => b:="2446";
                when 2447 => b:="2447";
                when 2448 => b:="2448";
                when 2449 => b:="2449";
                when 2450 => b:="2450";
                when 2451 => b:="2451";
                when 2452 => b:="2452";
                when 2453 => b:="2453";
                when 2454 => b:="2454";
                when 2455 => b:="2455";
                when 2456 => b:="2456";
                when 2457 => b:="2457";
                when 2458 => b:="2458";
                when 2459 => b:="2459";
                when 2460 => b:="2460";
                when 2461 => b:="2461";
                when 2462 => b:="2462";
                when 2463 => b:="2463";
                when 2464 => b:="2464";
                when 2465 => b:="2465";
                when 2466 => b:="2466";
                when 2467 => b:="2467";
                when 2468 => b:="2468";
                when 2469 => b:="2469";
                when 2470 => b:="2470";
                when 2471 => b:="2471";
                when 2472 => b:="2472";
                when 2473 => b:="2473";
                when 2474 => b:="2474";
                when 2475 => b:="2475";
                when 2476 => b:="2476";
                when 2477 => b:="2477";
                when 2478 => b:="2478";
                when 2479 => b:="2479";
                when 2480 => b:="2480";
                when 2481 => b:="2481";
                when 2482 => b:="2482";
                when 2483 => b:="2483";
                when 2484 => b:="2484";
                when 2485 => b:="2485";
                when 2486 => b:="2486";
                when 2487 => b:="2487";
                when 2488 => b:="2488";
                when 2489 => b:="2489";
                when 2490 => b:="2490";
                when 2491 => b:="2491";
                when 2492 => b:="2492";
                when 2493 => b:="2493";
                when 2494 => b:="2494";
                when 2495 => b:="2495";
                when 2496 => b:="2496";
                when 2497 => b:="2497";
                when 2498 => b:="2498";
                when 2499 => b:="2499";
                when 2500 => b:="2500";
                when 2501 => b:="2501";
                when 2502 => b:="2502";
                when 2503 => b:="2503";
                when 2504 => b:="2504";
                when 2505 => b:="2505";
                when 2506 => b:="2506";
                when 2507 => b:="2507";
                when 2508 => b:="2508";
                when 2509 => b:="2509";
                when 2510 => b:="2510";
                when 2511 => b:="2511";
                when 2512 => b:="2512";
                when 2513 => b:="2513";
                when 2514 => b:="2514";
                when 2515 => b:="2515";
                when 2516 => b:="2516";
                when 2517 => b:="2517";
                when 2518 => b:="2518";
                when 2519 => b:="2519";
                when 2520 => b:="2520";
                when 2521 => b:="2521";
                when 2522 => b:="2522";
                when 2523 => b:="2523";
                when 2524 => b:="2524";
                when 2525 => b:="2525";
                when 2526 => b:="2526";
                when 2527 => b:="2527";
                when 2528 => b:="2528";
                when 2529 => b:="2529";
                when 2530 => b:="2530";
                when 2531 => b:="2531";
                when 2532 => b:="2532";
                when 2533 => b:="2533";
                when 2534 => b:="2534";
                when 2535 => b:="2535";
                when 2536 => b:="2536";
                when 2537 => b:="2537";
                when 2538 => b:="2538";
                when 2539 => b:="2539";
                when 2540 => b:="2540";
                when 2541 => b:="2541";
                when 2542 => b:="2542";
                when 2543 => b:="2543";
                when 2544 => b:="2544";
                when 2545 => b:="2545";
                when 2546 => b:="2546";
                when 2547 => b:="2547";
                when 2548 => b:="2548";
                when 2549 => b:="2549";
                when 2550 => b:="2550";
                when 2551 => b:="2551";
                when 2552 => b:="2552";
                when 2553 => b:="2553";
                when 2554 => b:="2554";
                when 2555 => b:="2555";
                when 2556 => b:="2556";
                when 2557 => b:="2557";
                when 2558 => b:="2558";
                when 2559 => b:="2559";
                when 2560 => b:="2560";
                when 2561 => b:="2561";
                when 2562 => b:="2562";
                when 2563 => b:="2563";
                when 2564 => b:="2564";
                when 2565 => b:="2565";
                when 2566 => b:="2566";
                when 2567 => b:="2567";
                when 2568 => b:="2568";
                when 2569 => b:="2569";
                when 2570 => b:="2570";
                when 2571 => b:="2571";
                when 2572 => b:="2572";
                when 2573 => b:="2573";
                when 2574 => b:="2574";
                when 2575 => b:="2575";
                when 2576 => b:="2576";
                when 2577 => b:="2577";
                when 2578 => b:="2578";
                when 2579 => b:="2579";
                when 2580 => b:="2580";
                when 2581 => b:="2581";
                when 2582 => b:="2582";
                when 2583 => b:="2583";
                when 2584 => b:="2584";
                when 2585 => b:="2585";
                when 2586 => b:="2586";
                when 2587 => b:="2587";
                when 2588 => b:="2588";
                when 2589 => b:="2589";
                when 2590 => b:="2590";
                when 2591 => b:="2591";
                when 2592 => b:="2592";
                when 2593 => b:="2593";
                when 2594 => b:="2594";
                when 2595 => b:="2595";
                when 2596 => b:="2596";
                when 2597 => b:="2597";
                when 2598 => b:="2598";
                when 2599 => b:="2599";
                when 2600 => b:="2600";
                when 2601 => b:="2601";
                when 2602 => b:="2602";
                when 2603 => b:="2603";
                when 2604 => b:="2604";
                when 2605 => b:="2605";
                when 2606 => b:="2606";
                when 2607 => b:="2607";
                when 2608 => b:="2608";
                when 2609 => b:="2609";
                when 2610 => b:="2610";
                when 2611 => b:="2611";
                when 2612 => b:="2612";
                when 2613 => b:="2613";
                when 2614 => b:="2614";
                when 2615 => b:="2615";
                when 2616 => b:="2616";
                when 2617 => b:="2617";
                when 2618 => b:="2618";
                when 2619 => b:="2619";
                when 2620 => b:="2620";
                when 2621 => b:="2621";
                when 2622 => b:="2622";
                when 2623 => b:="2623";
                when 2624 => b:="2624";
                when 2625 => b:="2625";
                when 2626 => b:="2626";
                when 2627 => b:="2627";
                when 2628 => b:="2628";
                when 2629 => b:="2629";
                when 2630 => b:="2630";
                when 2631 => b:="2631";
                when 2632 => b:="2632";
                when 2633 => b:="2633";
                when 2634 => b:="2634";
                when 2635 => b:="2635";
                when 2636 => b:="2636";
                when 2637 => b:="2637";
                when 2638 => b:="2638";
                when 2639 => b:="2639";
                when 2640 => b:="2640";
                when 2641 => b:="2641";
                when 2642 => b:="2642";
                when 2643 => b:="2643";
                when 2644 => b:="2644";
                when 2645 => b:="2645";
                when 2646 => b:="2646";
                when 2647 => b:="2647";
                when 2648 => b:="2648";
                when 2649 => b:="2649";
                when 2650 => b:="2650";
                when 2651 => b:="2651";
                when 2652 => b:="2652";
                when 2653 => b:="2653";
                when 2654 => b:="2654";
                when 2655 => b:="2655";
                when 2656 => b:="2656";
                when 2657 => b:="2657";
                when 2658 => b:="2658";
                when 2659 => b:="2659";
                when 2660 => b:="2660";
                when 2661 => b:="2661";
                when 2662 => b:="2662";
                when 2663 => b:="2663";
                when 2664 => b:="2664";
                when 2665 => b:="2665";
                when 2666 => b:="2666";
                when 2667 => b:="2667";
                when 2668 => b:="2668";
                when 2669 => b:="2669";
                when 2670 => b:="2670";
                when 2671 => b:="2671";
                when 2672 => b:="2672";
                when 2673 => b:="2673";
                when 2674 => b:="2674";
                when 2675 => b:="2675";
                when 2676 => b:="2676";
                when 2677 => b:="2677";
                when 2678 => b:="2678";
                when 2679 => b:="2679";
                when 2680 => b:="2680";
                when 2681 => b:="2681";
                when 2682 => b:="2682";
                when 2683 => b:="2683";
                when 2684 => b:="2684";
                when 2685 => b:="2685";
                when 2686 => b:="2686";
                when 2687 => b:="2687";
                when 2688 => b:="2688";
                when 2689 => b:="2689";
                when 2690 => b:="2690";
                when 2691 => b:="2691";
                when 2692 => b:="2692";
                when 2693 => b:="2693";
                when 2694 => b:="2694";
                when 2695 => b:="2695";
                when 2696 => b:="2696";
                when 2697 => b:="2697";
                when 2698 => b:="2698";
                when 2699 => b:="2699";
                when 2700 => b:="2700";
                when 2701 => b:="2701";
                when 2702 => b:="2702";
                when 2703 => b:="2703";
                when 2704 => b:="2704";
                when 2705 => b:="2705";
                when 2706 => b:="2706";
                when 2707 => b:="2707";
                when 2708 => b:="2708";
                when 2709 => b:="2709";
                when 2710 => b:="2710";
                when 2711 => b:="2711";
                when 2712 => b:="2712";
                when 2713 => b:="2713";
                when 2714 => b:="2714";
                when 2715 => b:="2715";
                when 2716 => b:="2716";
                when 2717 => b:="2717";
                when 2718 => b:="2718";
                when 2719 => b:="2719";
                when 2720 => b:="2720";
                when 2721 => b:="2721";
                when 2722 => b:="2722";
                when 2723 => b:="2723";
                when 2724 => b:="2724";
                when 2725 => b:="2725";
                when 2726 => b:="2726";
                when 2727 => b:="2727";
                when 2728 => b:="2728";
                when 2729 => b:="2729";
                when 2730 => b:="2730";
                when 2731 => b:="2731";
                when 2732 => b:="2732";
                when 2733 => b:="2733";
                when 2734 => b:="2734";
                when 2735 => b:="2735";
                when 2736 => b:="2736";
                when 2737 => b:="2737";
                when 2738 => b:="2738";
                when 2739 => b:="2739";
                when 2740 => b:="2740";
                when 2741 => b:="2741";
                when 2742 => b:="2742";
                when 2743 => b:="2743";
                when 2744 => b:="2744";
                when 2745 => b:="2745";
                when 2746 => b:="2746";
                when 2747 => b:="2747";
                when 2748 => b:="2748";
                when 2749 => b:="2749";
                when 2750 => b:="2750";
                when 2751 => b:="2751";
                when 2752 => b:="2752";
                when 2753 => b:="2753";
                when 2754 => b:="2754";
                when 2755 => b:="2755";
                when 2756 => b:="2756";
                when 2757 => b:="2757";
                when 2758 => b:="2758";
                when 2759 => b:="2759";
                when 2760 => b:="2760";
                when 2761 => b:="2761";
                when 2762 => b:="2762";
                when 2763 => b:="2763";
                when 2764 => b:="2764";
                when 2765 => b:="2765";
                when 2766 => b:="2766";
                when 2767 => b:="2767";
                when 2768 => b:="2768";
                when 2769 => b:="2769";
                when 2770 => b:="2770";
                when 2771 => b:="2771";
                when 2772 => b:="2772";
                when 2773 => b:="2773";
                when 2774 => b:="2774";
                when 2775 => b:="2775";
                when 2776 => b:="2776";
                when 2777 => b:="2777";
                when 2778 => b:="2778";
                when 2779 => b:="2779";
                when 2780 => b:="2780";
                when 2781 => b:="2781";
                when 2782 => b:="2782";
                when 2783 => b:="2783";
                when 2784 => b:="2784";
                when 2785 => b:="2785";
                when 2786 => b:="2786";
                when 2787 => b:="2787";
                when 2788 => b:="2788";
                when 2789 => b:="2789";
                when 2790 => b:="2790";
                when 2791 => b:="2791";
                when 2792 => b:="2792";
                when 2793 => b:="2793";
                when 2794 => b:="2794";
                when 2795 => b:="2795";
                when 2796 => b:="2796";
                when 2797 => b:="2797";
                when 2798 => b:="2798";
                when 2799 => b:="2799";
                when 2800 => b:="2800";
                when 2801 => b:="2801";
                when 2802 => b:="2802";
                when 2803 => b:="2803";
                when 2804 => b:="2804";
                when 2805 => b:="2805";
                when 2806 => b:="2806";
                when 2807 => b:="2807";
                when 2808 => b:="2808";
                when 2809 => b:="2809";
                when 2810 => b:="2810";
                when 2811 => b:="2811";
                when 2812 => b:="2812";
                when 2813 => b:="2813";
                when 2814 => b:="2814";
                when 2815 => b:="2815";
                when 2816 => b:="2816";
                when 2817 => b:="2817";
                when 2818 => b:="2818";
                when 2819 => b:="2819";
                when 2820 => b:="2820";
                when 2821 => b:="2821";
                when 2822 => b:="2822";
                when 2823 => b:="2823";
                when 2824 => b:="2824";
                when 2825 => b:="2825";
                when 2826 => b:="2826";
                when 2827 => b:="2827";
                when 2828 => b:="2828";
                when 2829 => b:="2829";
                when 2830 => b:="2830";
                when 2831 => b:="2831";
                when 2832 => b:="2832";
                when 2833 => b:="2833";
                when 2834 => b:="2834";
                when 2835 => b:="2835";
                when 2836 => b:="2836";
                when 2837 => b:="2837";
                when 2838 => b:="2838";
                when 2839 => b:="2839";
                when 2840 => b:="2840";
                when 2841 => b:="2841";
                when 2842 => b:="2842";
                when 2843 => b:="2843";
                when 2844 => b:="2844";
                when 2845 => b:="2845";
                when 2846 => b:="2846";
                when 2847 => b:="2847";
                when 2848 => b:="2848";
                when 2849 => b:="2849";
                when 2850 => b:="2850";
                when 2851 => b:="2851";
                when 2852 => b:="2852";
                when 2853 => b:="2853";
                when 2854 => b:="2854";
                when 2855 => b:="2855";
                when 2856 => b:="2856";
                when 2857 => b:="2857";
                when 2858 => b:="2858";
                when 2859 => b:="2859";
                when 2860 => b:="2860";
                when 2861 => b:="2861";
                when 2862 => b:="2862";
                when 2863 => b:="2863";
                when 2864 => b:="2864";
                when 2865 => b:="2865";
                when 2866 => b:="2866";
                when 2867 => b:="2867";
                when 2868 => b:="2868";
                when 2869 => b:="2869";
                when 2870 => b:="2870";
                when 2871 => b:="2871";
                when 2872 => b:="2872";
                when 2873 => b:="2873";
                when 2874 => b:="2874";
                when 2875 => b:="2875";
                when 2876 => b:="2876";
                when 2877 => b:="2877";
                when 2878 => b:="2878";
                when 2879 => b:="2879";
                when 2880 => b:="2880";
                when 2881 => b:="2881";
                when 2882 => b:="2882";
                when 2883 => b:="2883";
                when 2884 => b:="2884";
                when 2885 => b:="2885";
                when 2886 => b:="2886";
                when 2887 => b:="2887";
                when 2888 => b:="2888";
                when 2889 => b:="2889";
                when 2890 => b:="2890";
                when 2891 => b:="2891";
                when 2892 => b:="2892";
                when 2893 => b:="2893";
                when 2894 => b:="2894";
                when 2895 => b:="2895";
                when 2896 => b:="2896";
                when 2897 => b:="2897";
                when 2898 => b:="2898";
                when 2899 => b:="2899";
                when 2900 => b:="2900";
                when 2901 => b:="2901";
                when 2902 => b:="2902";
                when 2903 => b:="2903";
                when 2904 => b:="2904";
                when 2905 => b:="2905";
                when 2906 => b:="2906";
                when 2907 => b:="2907";
                when 2908 => b:="2908";
                when 2909 => b:="2909";
                when 2910 => b:="2910";
                when 2911 => b:="2911";
                when 2912 => b:="2912";
                when 2913 => b:="2913";
                when 2914 => b:="2914";
                when 2915 => b:="2915";
                when 2916 => b:="2916";
                when 2917 => b:="2917";
                when 2918 => b:="2918";
                when 2919 => b:="2919";
                when 2920 => b:="2920";
                when 2921 => b:="2921";
                when 2922 => b:="2922";
                when 2923 => b:="2923";
                when 2924 => b:="2924";
                when 2925 => b:="2925";
                when 2926 => b:="2926";
                when 2927 => b:="2927";
                when 2928 => b:="2928";
                when 2929 => b:="2929";
                when 2930 => b:="2930";
                when 2931 => b:="2931";
                when 2932 => b:="2932";
                when 2933 => b:="2933";
                when 2934 => b:="2934";
                when 2935 => b:="2935";
                when 2936 => b:="2936";
                when 2937 => b:="2937";
                when 2938 => b:="2938";
                when 2939 => b:="2939";
                when 2940 => b:="2940";
                when 2941 => b:="2941";
                when 2942 => b:="2942";
                when 2943 => b:="2943";
                when 2944 => b:="2944";
                when 2945 => b:="2945";
                when 2946 => b:="2946";
                when 2947 => b:="2947";
                when 2948 => b:="2948";
                when 2949 => b:="2949";
                when 2950 => b:="2950";
                when 2951 => b:="2951";
                when 2952 => b:="2952";
                when 2953 => b:="2953";
                when 2954 => b:="2954";
                when 2955 => b:="2955";
                when 2956 => b:="2956";
                when 2957 => b:="2957";
                when 2958 => b:="2958";
                when 2959 => b:="2959";
                when 2960 => b:="2960";
                when 2961 => b:="2961";
                when 2962 => b:="2962";
                when 2963 => b:="2963";
                when 2964 => b:="2964";
                when 2965 => b:="2965";
                when 2966 => b:="2966";
                when 2967 => b:="2967";
                when 2968 => b:="2968";
                when 2969 => b:="2969";
                when 2970 => b:="2970";
                when 2971 => b:="2971";
                when 2972 => b:="2972";
                when 2973 => b:="2973";
                when 2974 => b:="2974";
                when 2975 => b:="2975";
                when 2976 => b:="2976";
                when 2977 => b:="2977";
                when 2978 => b:="2978";
                when 2979 => b:="2979";
                when 2980 => b:="2980";
                when 2981 => b:="2981";
                when 2982 => b:="2982";
                when 2983 => b:="2983";
                when 2984 => b:="2984";
                when 2985 => b:="2985";
                when 2986 => b:="2986";
                when 2987 => b:="2987";
                when 2988 => b:="2988";
                when 2989 => b:="2989";
                when 2990 => b:="2990";
                when 2991 => b:="2991";
                when 2992 => b:="2992";
                when 2993 => b:="2993";
                when 2994 => b:="2994";
                when 2995 => b:="2995";
                when 2996 => b:="2996";
                when 2997 => b:="2997";
                when 2998 => b:="2998";
                when 3000 => b:="3000";
                when 3001 => b:="3001";
                when 3002 => b:="3002";
                when 3003 => b:="3003";
                when 3004 => b:="3004";
                when 3005 => b:="3005";
                when 3006 => b:="3006";
                when 3007 => b:="3007";
                when 3008 => b:="3008";
                when 3009 => b:="3009";
                when 3010 => b:="3010";
                when 3011 => b:="3011";
                when 3012 => b:="3012";
                when 3013 => b:="3013";
                when 3014 => b:="3014";
                when 3015 => b:="3015";
                when 3016 => b:="3016";
                when 3017 => b:="3017";
                when 3018 => b:="3018";
                when 3019 => b:="3019";
                when 3020 => b:="3020";
                when 3021 => b:="3021";
                when 3022 => b:="3022";
                when 3023 => b:="3023";
                when 3024 => b:="3024";
                when 3025 => b:="3025";
                when 3026 => b:="3026";
                when 3027 => b:="3027";
                when 3028 => b:="3028";
                when 3029 => b:="3029";
                when 3030 => b:="3030";
                when 3031 => b:="3031";
                when 3032 => b:="3032";
                when 3033 => b:="3033";
                when 3034 => b:="3034";
                when 3035 => b:="3035";
                when 3036 => b:="3036";
                when 3037 => b:="3037";
                when 3038 => b:="3038";
                when 3039 => b:="3039";
                when 3040 => b:="3040";
                when 3041 => b:="3041";
                when 3042 => b:="3042";
                when 3043 => b:="3043";
                when 3044 => b:="3044";
                when 3045 => b:="3045";
                when 3046 => b:="3046";
                when 3047 => b:="3047";
                when 3048 => b:="3048";
                when 3049 => b:="3049";
                when 3050 => b:="3050";
                when 3051 => b:="3051";
                when 3052 => b:="3052";
                when 3053 => b:="3053";
                when 3054 => b:="3054";
                when 3055 => b:="3055";
                when 3056 => b:="3056";
                when 3057 => b:="3057";
                when 3058 => b:="3058";
                when 3059 => b:="3059";
                when 3060 => b:="3060";
                when 3061 => b:="3061";
                when 3062 => b:="3062";
                when 3063 => b:="3063";
                when 3064 => b:="3064";
                when 3065 => b:="3065";
                when 3066 => b:="3066";
                when 3067 => b:="3067";
                when 3068 => b:="3068";
                when 3069 => b:="3069";
                when 3070 => b:="3070";
                when 3071 => b:="3071";
                when 3072 => b:="3072";
                when 3073 => b:="3073";
                when 3074 => b:="3074";
                when 3075 => b:="3075";
                when 3076 => b:="3076";
                when 3077 => b:="3077";
                when 3078 => b:="3078";
                when 3079 => b:="3079";
                when 3080 => b:="3080";
                when 3081 => b:="3081";
                when 3082 => b:="3082";
                when 3083 => b:="3083";
                when 3084 => b:="3084";
                when 3085 => b:="3085";
                when 3086 => b:="3086";
                when 3087 => b:="3087";
                when 3088 => b:="3088";
                when 3089 => b:="3089";
                when 3090 => b:="3090";
                when 3091 => b:="3091";
                when 3092 => b:="3092";
                when 3093 => b:="3093";
                when 3094 => b:="3094";
                when 3095 => b:="3095";
                when 3096 => b:="3096";
                when 3097 => b:="3097";
                when 3098 => b:="3098";
                when 3099 => b:="3099";
                when 3100 => b:="3100";
                when 3101 => b:="3101";
                when 3102 => b:="3102";
                when 3103 => b:="3103";
                when 3104 => b:="3104";
                when 3105 => b:="3105";
                when 3106 => b:="3106";
                when 3107 => b:="3107";
                when 3108 => b:="3108";
                when 3109 => b:="3109";
                when 3110 => b:="3110";
                when 3111 => b:="3111";
                when 3112 => b:="3112";
                when 3113 => b:="3113";
                when 3114 => b:="3114";
                when 3115 => b:="3115";
                when 3116 => b:="3116";
                when 3117 => b:="3117";
                when 3118 => b:="3118";
                when 3119 => b:="3119";
                when 3120 => b:="3120";
                when 3121 => b:="3121";
                when 3122 => b:="3122";
                when 3123 => b:="3123";
                when 3124 => b:="3124";
                when 3125 => b:="3125";
                when 3126 => b:="3126";
                when 3127 => b:="3127";
                when 3128 => b:="3128";
                when 3129 => b:="3129";
                when 3130 => b:="3130";
                when 3131 => b:="3131";
                when 3132 => b:="3132";
                when 3133 => b:="3133";
                when 3134 => b:="3134";
                when 3135 => b:="3135";
                when 3136 => b:="3136";
                when 3137 => b:="3137";
                when 3138 => b:="3138";
                when 3139 => b:="3139";
                when 3140 => b:="3140";
                when 3141 => b:="3141";
                when 3142 => b:="3142";
                when 3143 => b:="3143";
                when 3144 => b:="3144";
                when 3145 => b:="3145";
                when 3146 => b:="3146";
                when 3147 => b:="3147";
                when 3148 => b:="3148";
                when 3149 => b:="3149";
                when 3150 => b:="3150";
                when 3151 => b:="3151";
                when 3152 => b:="3152";
                when 3153 => b:="3153";
                when 3154 => b:="3154";
                when 3155 => b:="3155";
                when 3156 => b:="3156";
                when 3157 => b:="3157";
                when 3158 => b:="3158";
                when 3159 => b:="3159";
                when 3160 => b:="3160";
                when 3161 => b:="3161";
                when 3162 => b:="3162";
                when 3163 => b:="3163";
                when 3164 => b:="3164";
                when 3165 => b:="3165";
                when 3166 => b:="3166";
                when 3167 => b:="3167";
                when 3168 => b:="3168";
                when 3169 => b:="3169";
                when 3170 => b:="3170";
                when 3171 => b:="3171";
                when 3172 => b:="3172";
                when 3173 => b:="3173";
                when 3174 => b:="3174";
                when 3175 => b:="3175";
                when 3176 => b:="3176";
                when 3177 => b:="3177";
                when 3178 => b:="3178";
                when 3179 => b:="3179";
                when 3180 => b:="3180";
                when 3181 => b:="3181";
                when 3182 => b:="3182";
                when 3183 => b:="3183";
                when 3184 => b:="3184";
                when 3185 => b:="3185";
                when 3186 => b:="3186";
                when 3187 => b:="3187";
                when 3188 => b:="3188";
                when 3189 => b:="3189";
                when 3190 => b:="3190";
                when 3191 => b:="3191";
                when 3192 => b:="3192";
                when 3193 => b:="3193";
                when 3194 => b:="3194";
                when 3195 => b:="3195";
                when 3196 => b:="3196";
                when 3197 => b:="3197";
                when 3198 => b:="3198";
                when 3199 => b:="3199";
                when 3200 => b:="3200";
                when 3201 => b:="3201";
                when 3202 => b:="3202";
                when 3203 => b:="3203";
                when 3204 => b:="3204";
                when 3205 => b:="3205";
                when 3206 => b:="3206";
                when 3207 => b:="3207";
                when 3208 => b:="3208";
                when 3209 => b:="3209";
                when 3210 => b:="3210";
                when 3211 => b:="3211";
                when 3212 => b:="3212";
                when 3213 => b:="3213";
                when 3214 => b:="3214";
                when 3215 => b:="3215";
                when 3216 => b:="3216";
                when 3217 => b:="3217";
                when 3218 => b:="3218";
                when 3219 => b:="3219";
                when 3220 => b:="3220";
                when 3221 => b:="3221";
                when 3222 => b:="3222";
                when 3223 => b:="3223";
                when 3224 => b:="3224";
                when 3225 => b:="3225";
                when 3226 => b:="3226";
                when 3227 => b:="3227";
                when 3228 => b:="3228";
                when 3229 => b:="3229";
                when 3230 => b:="3230";
                when 3231 => b:="3231";
                when 3232 => b:="3232";
                when 3233 => b:="3233";
                when 3234 => b:="3234";
                when 3235 => b:="3235";
                when 3236 => b:="3236";
                when 3237 => b:="3237";
                when 3238 => b:="3238";
                when 3239 => b:="3239";
                when 3240 => b:="3240";
                when 3241 => b:="3241";
                when 3242 => b:="3242";
                when 3243 => b:="3243";
                when 3244 => b:="3244";
                when 3245 => b:="3245";
                when 3246 => b:="3246";
                when 3247 => b:="3247";
                when 3248 => b:="3248";
                when 3249 => b:="3249";
                when 3250 => b:="3250";
                when 3251 => b:="3251";
                when 3252 => b:="3252";
                when 3253 => b:="3253";
                when 3254 => b:="3254";
                when 3255 => b:="3255";
                when 3256 => b:="3256";
                when 3257 => b:="3257";
                when 3258 => b:="3258";
                when 3259 => b:="3259";
                when 3260 => b:="3260";
                when 3261 => b:="3261";
                when 3262 => b:="3262";
                when 3263 => b:="3263";
                when 3264 => b:="3264";
                when 3265 => b:="3265";
                when 3266 => b:="3266";
                when 3267 => b:="3267";
                when 3268 => b:="3268";
                when 3269 => b:="3269";
                when 3270 => b:="3270";
                when 3271 => b:="3271";
                when 3272 => b:="3272";
                when 3273 => b:="3273";
                when 3274 => b:="3274";
                when 3275 => b:="3275";
                when 3276 => b:="3276";
                when 3277 => b:="3277";
                when 3278 => b:="3278";
                when 3279 => b:="3279";
                when 3280 => b:="3280";
                when 3281 => b:="3281";
                when 3282 => b:="3282";
                when 3283 => b:="3283";
                when 3284 => b:="3284";
                when 3285 => b:="3285";
                when 3286 => b:="3286";
                when 3287 => b:="3287";
                when 3288 => b:="3288";
                when 3289 => b:="3289";
                when 3290 => b:="3290";
                when 3291 => b:="3291";
                when 3292 => b:="3292";
                when 3293 => b:="3293";
                when 3294 => b:="3294";
                when 3295 => b:="3295";
                when 3296 => b:="3296";
                when 3297 => b:="3297";
                when 3298 => b:="3298";
                when 3299 => b:="3299";
                when 3300 => b:="3300";
                when 3301 => b:="3301";
                when 3302 => b:="3302";
                when 3303 => b:="3303";
                when 3304 => b:="3304";
                when 3305 => b:="3305";
                when 3306 => b:="3306";
                when 3307 => b:="3307";
                when 3308 => b:="3308";
                when 3309 => b:="3309";
                when 3310 => b:="3310";
                when 3311 => b:="3311";
                when 3312 => b:="3312";
                when 3313 => b:="3313";
                when 3314 => b:="3314";
                when 3315 => b:="3315";
                when 3316 => b:="3316";
                when 3317 => b:="3317";
                when 3318 => b:="3318";
                when 3319 => b:="3319";
                when 3320 => b:="3320";
                when 3321 => b:="3321";
                when 3322 => b:="3322";
                when 3323 => b:="3323";
                when 3324 => b:="3324";
                when 3325 => b:="3325";
                when 3326 => b:="3326";
                when 3327 => b:="3327";
                when 3328 => b:="3328";
                when 3329 => b:="3329";
                when 3330 => b:="3330";
                when 3331 => b:="3331";
                when 3332 => b:="3332";
                when 3333 => b:="3333";
                when 3334 => b:="3334";
                when 3335 => b:="3335";
                when 3336 => b:="3336";
                when 3337 => b:="3337";
                when 3338 => b:="3338";
                when 3339 => b:="3339";
                when 3340 => b:="3340";
                when 3341 => b:="3341";
                when 3342 => b:="3342";
                when 3343 => b:="3343";
                when 3344 => b:="3344";
                when 3345 => b:="3345";
                when 3346 => b:="3346";
                when 3347 => b:="3347";
                when 3348 => b:="3348";
                when 3349 => b:="3349";
                when 3350 => b:="3350";
                when 3351 => b:="3351";
                when 3352 => b:="3352";
                when 3353 => b:="3353";
                when 3354 => b:="3354";
                when 3355 => b:="3355";
                when 3356 => b:="3356";
                when 3357 => b:="3357";
                when 3358 => b:="3358";
                when 3359 => b:="3359";
                when 3360 => b:="3360";
                when 3361 => b:="3361";
                when 3362 => b:="3362";
                when 3363 => b:="3363";
                when 3364 => b:="3364";
                when 3365 => b:="3365";
                when 3366 => b:="3366";
                when 3367 => b:="3367";
                when 3368 => b:="3368";
                when 3369 => b:="3369";
                when 3370 => b:="3370";
                when 3371 => b:="3371";
                when 3372 => b:="3372";
                when 3373 => b:="3373";
                when 3374 => b:="3374";
                when 3375 => b:="3375";
                when 3376 => b:="3376";
                when 3377 => b:="3377";
                when 3378 => b:="3378";
                when 3379 => b:="3379";
                when 3380 => b:="3380";
                when 3381 => b:="3381";
                when 3382 => b:="3382";
                when 3383 => b:="3383";
                when 3384 => b:="3384";
                when 3385 => b:="3385";
                when 3386 => b:="3386";
                when 3387 => b:="3387";
                when 3388 => b:="3388";
                when 3389 => b:="3389";
                when 3390 => b:="3390";
                when 3391 => b:="3391";
                when 3392 => b:="3392";
                when 3393 => b:="3393";
                when 3394 => b:="3394";
                when 3395 => b:="3395";
                when 3396 => b:="3396";
                when 3397 => b:="3397";
                when 3398 => b:="3398";
                when 3399 => b:="3399";
                when 3400 => b:="3400";
                when 3401 => b:="3401";
                when 3402 => b:="3402";
                when 3403 => b:="3403";
                when 3404 => b:="3404";
                when 3405 => b:="3405";
                when 3406 => b:="3406";
                when 3407 => b:="3407";
                when 3408 => b:="3408";
                when 3409 => b:="3409";
                when 3410 => b:="3410";
                when 3411 => b:="3411";
                when 3412 => b:="3412";
                when 3413 => b:="3413";
                when 3414 => b:="3414";
                when 3415 => b:="3415";
                when 3416 => b:="3416";
                when 3417 => b:="3417";
                when 3418 => b:="3418";
                when 3419 => b:="3419";
                when 3420 => b:="3420";
                when 3421 => b:="3421";
                when 3422 => b:="3422";
                when 3423 => b:="3423";
                when 3424 => b:="3424";
                when 3425 => b:="3425";
                when 3426 => b:="3426";
                when 3427 => b:="3427";
                when 3428 => b:="3428";
                when 3429 => b:="3429";
                when 3430 => b:="3430";
                when 3431 => b:="3431";
                when 3432 => b:="3432";
                when 3433 => b:="3433";
                when 3434 => b:="3434";
                when 3435 => b:="3435";
                when 3436 => b:="3436";
                when 3437 => b:="3437";
                when 3438 => b:="3438";
                when 3439 => b:="3439";
                when 3440 => b:="3440";
                when 3441 => b:="3441";
                when 3442 => b:="3442";
                when 3443 => b:="3443";
                when 3444 => b:="3444";
                when 3445 => b:="3445";
                when 3446 => b:="3446";
                when 3447 => b:="3447";
                when 3448 => b:="3448";
                when 3449 => b:="3449";
                when 3450 => b:="3450";
                when 3451 => b:="3451";
                when 3452 => b:="3452";
                when 3453 => b:="3453";
                when 3454 => b:="3454";
                when 3455 => b:="3455";
                when 3456 => b:="3456";
                when 3457 => b:="3457";
                when 3458 => b:="3458";
                when 3459 => b:="3459";
                when 3460 => b:="3460";
                when 3461 => b:="3461";
                when 3462 => b:="3462";
                when 3463 => b:="3463";
                when 3464 => b:="3464";
                when 3465 => b:="3465";
                when 3466 => b:="3466";
                when 3467 => b:="3467";
                when 3468 => b:="3468";
                when 3469 => b:="3469";
                when 3470 => b:="3470";
                when 3471 => b:="3471";
                when 3472 => b:="3472";
                when 3473 => b:="3473";
                when 3474 => b:="3474";
                when 3475 => b:="3475";
                when 3476 => b:="3476";
                when 3477 => b:="3477";
                when 3478 => b:="3478";
                when 3479 => b:="3479";
                when 3480 => b:="3480";
                when 3481 => b:="3481";
                when 3482 => b:="3482";
                when 3483 => b:="3483";
                when 3484 => b:="3484";
                when 3485 => b:="3485";
                when 3486 => b:="3486";
                when 3487 => b:="3487";
                when 3488 => b:="3488";
                when 3489 => b:="3489";
                when 3490 => b:="3490";
                when 3491 => b:="3491";
                when 3492 => b:="3492";
                when 3493 => b:="3493";
                when 3494 => b:="3494";
                when 3495 => b:="3495";
                when 3496 => b:="3496";
                when 3497 => b:="3497";
                when 3498 => b:="3498";
                when 3499 => b:="3499";
                when 3500 => b:="3500";
                when 3501 => b:="3501";
                when 3502 => b:="3502";
                when 3503 => b:="3503";
                when 3504 => b:="3504";
                when 3505 => b:="3505";
                when 3506 => b:="3506";
                when 3507 => b:="3507";
                when 3508 => b:="3508";
                when 3509 => b:="3509";
                when 3510 => b:="3510";
                when 3511 => b:="3511";
                when 3512 => b:="3512";
                when 3513 => b:="3513";
                when 3514 => b:="3514";
                when 3515 => b:="3515";
                when 3516 => b:="3516";
                when 3517 => b:="3517";
                when 3518 => b:="3518";
                when 3519 => b:="3519";
                when 3520 => b:="3520";
                when 3521 => b:="3521";
                when 3522 => b:="3522";
                when 3523 => b:="3523";
                when 3524 => b:="3524";
                when 3525 => b:="3525";
                when 3526 => b:="3526";
                when 3527 => b:="3527";
                when 3528 => b:="3528";
                when 3529 => b:="3529";
                when 3530 => b:="3530";
                when 3531 => b:="3531";
                when 3532 => b:="3532";
                when 3533 => b:="3533";
                when 3534 => b:="3534";
                when 3535 => b:="3535";
                when 3536 => b:="3536";
                when 3537 => b:="3537";
                when 3538 => b:="3538";
                when 3539 => b:="3539";
                when 3540 => b:="3540";
                when 3541 => b:="3541";
                when 3542 => b:="3542";
                when 3543 => b:="3543";
                when 3544 => b:="3544";
                when 3545 => b:="3545";
                when 3546 => b:="3546";
                when 3547 => b:="3547";
                when 3548 => b:="3548";
                when 3549 => b:="3549";
                when 3550 => b:="3550";
                when 3551 => b:="3551";
                when 3552 => b:="3552";
                when 3553 => b:="3553";
                when 3554 => b:="3554";
                when 3555 => b:="3555";
                when 3556 => b:="3556";
                when 3557 => b:="3557";
                when 3558 => b:="3558";
                when 3559 => b:="3559";
                when 3560 => b:="3560";
                when 3561 => b:="3561";
                when 3562 => b:="3562";
                when 3563 => b:="3563";
                when 3564 => b:="3564";
                when 3565 => b:="3565";
                when 3566 => b:="3566";
                when 3567 => b:="3567";
                when 3568 => b:="3568";
                when 3569 => b:="3569";
                when 3570 => b:="3570";
                when 3571 => b:="3571";
                when 3572 => b:="3572";
                when 3573 => b:="3573";
                when 3574 => b:="3574";
                when 3575 => b:="3575";
                when 3576 => b:="3576";
                when 3577 => b:="3577";
                when 3578 => b:="3578";
                when 3579 => b:="3579";
                when 3580 => b:="3580";
                when 3581 => b:="3581";
                when 3582 => b:="3582";
                when 3583 => b:="3583";
                when 3584 => b:="3584";
                when 3585 => b:="3585";
                when 3586 => b:="3586";
                when 3587 => b:="3587";
                when 3588 => b:="3588";
                when 3589 => b:="3589";
                when 3590 => b:="3590";
                when 3591 => b:="3591";
                when 3592 => b:="3592";
                when 3593 => b:="3593";
                when 3594 => b:="3594";
                when 3595 => b:="3595";
                when 3596 => b:="3596";
                when 3597 => b:="3597";
                when 3598 => b:="3598";
                when 3599 => b:="3599";
                when 3600 => b:="3600";
                when 3601 => b:="3601";
                when 3602 => b:="3602";
                when 3603 => b:="3603";
                when 3604 => b:="3604";
                when 3605 => b:="3605";
                when 3606 => b:="3606";
                when 3607 => b:="3607";
                when 3608 => b:="3608";
                when 3609 => b:="3609";
                when 3610 => b:="3610";
                when 3611 => b:="3611";
                when 3612 => b:="3612";
                when 3613 => b:="3613";
                when 3614 => b:="3614";
                when 3615 => b:="3615";
                when 3616 => b:="3616";
                when 3617 => b:="3617";
                when 3618 => b:="3618";
                when 3619 => b:="3619";
                when 3620 => b:="3620";
                when 3621 => b:="3621";
                when 3622 => b:="3622";
                when 3623 => b:="3623";
                when 3624 => b:="3624";
                when 3625 => b:="3625";
                when 3626 => b:="3626";
                when 3627 => b:="3627";
                when 3628 => b:="3628";
                when 3629 => b:="3629";
                when 3630 => b:="3630";
                when 3631 => b:="3631";
                when 3632 => b:="3632";
                when 3633 => b:="3633";
                when 3634 => b:="3634";
                when 3635 => b:="3635";
                when 3636 => b:="3636";
                when 3637 => b:="3637";
                when 3638 => b:="3638";
                when 3639 => b:="3639";
                when 3640 => b:="3640";
                when 3641 => b:="3641";
                when 3642 => b:="3642";
                when 3643 => b:="3643";
                when 3644 => b:="3644";
                when 3645 => b:="3645";
                when 3646 => b:="3646";
                when 3647 => b:="3647";
                when 3648 => b:="3648";
                when 3649 => b:="3649";
                when 3650 => b:="3650";
                when 3651 => b:="3651";
                when 3652 => b:="3652";
                when 3653 => b:="3653";
                when 3654 => b:="3654";
                when 3655 => b:="3655";
                when 3656 => b:="3656";
                when 3657 => b:="3657";
                when 3658 => b:="3658";
                when 3659 => b:="3659";
                when 3660 => b:="3660";
                when 3661 => b:="3661";
                when 3662 => b:="3662";
                when 3663 => b:="3663";
                when 3664 => b:="3664";
                when 3665 => b:="3665";
                when 3666 => b:="3666";
                when 3667 => b:="3667";
                when 3668 => b:="3668";
                when 3669 => b:="3669";
                when 3670 => b:="3670";
                when 3671 => b:="3671";
                when 3672 => b:="3672";
                when 3673 => b:="3673";
                when 3674 => b:="3674";
                when 3675 => b:="3675";
                when 3676 => b:="3676";
                when 3677 => b:="3677";
                when 3678 => b:="3678";
                when 3679 => b:="3679";
                when 3680 => b:="3680";
                when 3681 => b:="3681";
                when 3682 => b:="3682";
                when 3683 => b:="3683";
                when 3684 => b:="3684";
                when 3685 => b:="3685";
                when 3686 => b:="3686";
                when 3687 => b:="3687";
                when 3688 => b:="3688";
                when 3689 => b:="3689";
                when 3690 => b:="3690";
                when 3691 => b:="3691";
                when 3692 => b:="3692";
                when 3693 => b:="3693";
                when 3694 => b:="3694";
                when 3695 => b:="3695";
                when 3696 => b:="3696";
                when 3697 => b:="3697";
                when 3698 => b:="3698";
                when 3699 => b:="3699";
                when 3700 => b:="3700";
                when 3701 => b:="3701";
                when 3702 => b:="3702";
                when 3703 => b:="3703";
                when 3704 => b:="3704";
                when 3705 => b:="3705";
                when 3706 => b:="3706";
                when 3707 => b:="3707";
                when 3708 => b:="3708";
                when 3709 => b:="3709";
                when 3710 => b:="3710";
                when 3711 => b:="3711";
                when 3712 => b:="3712";
                when 3713 => b:="3713";
                when 3714 => b:="3714";
                when 3715 => b:="3715";
                when 3716 => b:="3716";
                when 3717 => b:="3717";
                when 3718 => b:="3718";
                when 3719 => b:="3719";
                when 3720 => b:="3720";
                when 3721 => b:="3721";
                when 3722 => b:="3722";
                when 3723 => b:="3723";
                when 3724 => b:="3724";
                when 3725 => b:="3725";
                when 3726 => b:="3726";
                when 3727 => b:="3727";
                when 3728 => b:="3728";
                when 3729 => b:="3729";
                when 3730 => b:="3730";
                when 3731 => b:="3731";
                when 3732 => b:="3732";
                when 3733 => b:="3733";
                when 3734 => b:="3734";
                when 3735 => b:="3735";
                when 3736 => b:="3736";
                when 3737 => b:="3737";
                when 3738 => b:="3738";
                when 3739 => b:="3739";
                when 3740 => b:="3740";
                when 3741 => b:="3741";
                when 3742 => b:="3742";
                when 3743 => b:="3743";
                when 3744 => b:="3744";
                when 3745 => b:="3745";
                when 3746 => b:="3746";
                when 3747 => b:="3747";
                when 3748 => b:="3748";
                when 3749 => b:="3749";
                when 3750 => b:="3750";
                when 3751 => b:="3751";
                when 3752 => b:="3752";
                when 3753 => b:="3753";
                when 3754 => b:="3754";
                when 3755 => b:="3755";
                when 3756 => b:="3756";
                when 3757 => b:="3757";
                when 3758 => b:="3758";
                when 3759 => b:="3759";
                when 3760 => b:="3760";
                when 3761 => b:="3761";
                when 3762 => b:="3762";
                when 3763 => b:="3763";
                when 3764 => b:="3764";
                when 3765 => b:="3765";
                when 3766 => b:="3766";
                when 3767 => b:="3767";
                when 3768 => b:="3768";
                when 3769 => b:="3769";
                when 3770 => b:="3770";
                when 3771 => b:="3771";
                when 3772 => b:="3772";
                when 3773 => b:="3773";
                when 3774 => b:="3774";
                when 3775 => b:="3775";
                when 3776 => b:="3776";
                when 3777 => b:="3777";
                when 3778 => b:="3778";
                when 3779 => b:="3779";
                when 3780 => b:="3780";
                when 3781 => b:="3781";
                when 3782 => b:="3782";
                when 3783 => b:="3783";
                when 3784 => b:="3784";
                when 3785 => b:="3785";
                when 3786 => b:="3786";
                when 3787 => b:="3787";
                when 3788 => b:="3788";
                when 3789 => b:="3789";
                when 3790 => b:="3790";
                when 3791 => b:="3791";
                when 3792 => b:="3792";
                when 3793 => b:="3793";
                when 3794 => b:="3794";
                when 3795 => b:="3795";
                when 3796 => b:="3796";
                when 3797 => b:="3797";
                when 3798 => b:="3798";
                when 3799 => b:="3799";
                when 3800 => b:="3800";
                when 3801 => b:="3801";
                when 3802 => b:="3802";
                when 3803 => b:="3803";
                when 3804 => b:="3804";
                when 3805 => b:="3805";
                when 3806 => b:="3806";
                when 3807 => b:="3807";
                when 3808 => b:="3808";
                when 3809 => b:="3809";
                when 3810 => b:="3810";
                when 3811 => b:="3811";
                when 3812 => b:="3812";
                when 3813 => b:="3813";
                when 3814 => b:="3814";
                when 3815 => b:="3815";
                when 3816 => b:="3816";
                when 3817 => b:="3817";
                when 3818 => b:="3818";
                when 3819 => b:="3819";
                when 3820 => b:="3820";
                when 3821 => b:="3821";
                when 3822 => b:="3822";
                when 3823 => b:="3823";
                when 3824 => b:="3824";
                when 3825 => b:="3825";
                when 3826 => b:="3826";
                when 3827 => b:="3827";
                when 3828 => b:="3828";
                when 3829 => b:="3829";
                when 3830 => b:="3830";
                when 3831 => b:="3831";
                when 3832 => b:="3832";
                when 3833 => b:="3833";
                when 3834 => b:="3834";
                when 3835 => b:="3835";
                when 3836 => b:="3836";
                when 3837 => b:="3837";
                when 3838 => b:="3838";
                when 3839 => b:="3839";
                when 3840 => b:="3840";
                when 3841 => b:="3841";
                when 3842 => b:="3842";
                when 3843 => b:="3843";
                when 3844 => b:="3844";
                when 3845 => b:="3845";
                when 3846 => b:="3846";
                when 3847 => b:="3847";
                when 3848 => b:="3848";
                when 3849 => b:="3849";
                when 3850 => b:="3850";
                when 3851 => b:="3851";
                when 3852 => b:="3852";
                when 3853 => b:="3853";
                when 3854 => b:="3854";
                when 3855 => b:="3855";
                when 3856 => b:="3856";
                when 3857 => b:="3857";
                when 3858 => b:="3858";
                when 3859 => b:="3859";
                when 3860 => b:="3860";
                when 3861 => b:="3861";
                when 3862 => b:="3862";
                when 3863 => b:="3863";
                when 3864 => b:="3864";
                when 3865 => b:="3865";
                when 3866 => b:="3866";
                when 3867 => b:="3867";
                when 3868 => b:="3868";
                when 3869 => b:="3869";
                when 3870 => b:="3870";
                when 3871 => b:="3871";
                when 3872 => b:="3872";
                when 3873 => b:="3873";
                when 3874 => b:="3874";
                when 3875 => b:="3875";
                when 3876 => b:="3876";
                when 3877 => b:="3877";
                when 3878 => b:="3878";
                when 3879 => b:="3879";
                when 3880 => b:="3880";
                when 3881 => b:="3881";
                when 3882 => b:="3882";
                when 3883 => b:="3883";
                when 3884 => b:="3884";
                when 3885 => b:="3885";
                when 3886 => b:="3886";
                when 3887 => b:="3887";
                when 3888 => b:="3888";
                when 3889 => b:="3889";
                when 3890 => b:="3890";
                when 3891 => b:="3891";
                when 3892 => b:="3892";
                when 3893 => b:="3893";
                when 3894 => b:="3894";
                when 3895 => b:="3895";
                when 3896 => b:="3896";
                when 3897 => b:="3897";
                when 3898 => b:="3898";
                when 3899 => b:="3899";
                when 3900 => b:="3900";
                when 3901 => b:="3901";
                when 3902 => b:="3902";
                when 3903 => b:="3903";
                when 3904 => b:="3904";
                when 3905 => b:="3905";
                when 3906 => b:="3906";
                when 3907 => b:="3907";
                when 3908 => b:="3908";
                when 3909 => b:="3909";
                when 3910 => b:="3910";
                when 3911 => b:="3911";
                when 3912 => b:="3912";
                when 3913 => b:="3913";
                when 3914 => b:="3914";
                when 3915 => b:="3915";
                when 3916 => b:="3916";
                when 3917 => b:="3917";
                when 3918 => b:="3918";
                when 3919 => b:="3919";
                when 3920 => b:="3920";
                when 3921 => b:="3921";
                when 3922 => b:="3922";
                when 3923 => b:="3923";
                when 3924 => b:="3924";
                when 3925 => b:="3925";
                when 3926 => b:="3926";
                when 3927 => b:="3927";
                when 3928 => b:="3928";
                when 3929 => b:="3929";
                when 3930 => b:="3930";
                when 3931 => b:="3931";
                when 3932 => b:="3932";
                when 3933 => b:="3933";
                when 3934 => b:="3934";
                when 3935 => b:="3935";
                when 3936 => b:="3936";
                when 3937 => b:="3937";
                when 3938 => b:="3938";
                when 3939 => b:="3939";
                when 3940 => b:="3940";
                when 3941 => b:="3941";
                when 3942 => b:="3942";
                when 3943 => b:="3943";
                when 3944 => b:="3944";
                when 3945 => b:="3945";
                when 3946 => b:="3946";
                when 3947 => b:="3947";
                when 3948 => b:="3948";
                when 3949 => b:="3949";
                when 3950 => b:="3950";
                when 3951 => b:="3951";
                when 3952 => b:="3952";
                when 3953 => b:="3953";
                when 3954 => b:="3954";
                when 3955 => b:="3955";
                when 3956 => b:="3956";
                when 3957 => b:="3957";
                when 3958 => b:="3958";
                when 3959 => b:="3959";
                when 3960 => b:="3960";
                when 3961 => b:="3961";
                when 3962 => b:="3962";
                when 3963 => b:="3963";
                when 3964 => b:="3964";
                when 3965 => b:="3965";
                when 3966 => b:="3966";
                when 3967 => b:="3967";
                when 3968 => b:="3968";
                when 3969 => b:="3969";
                when 3970 => b:="3970";
                when 3971 => b:="3971";
                when 3972 => b:="3972";
                when 3973 => b:="3973";
                when 3974 => b:="3974";
                when 3975 => b:="3975";
                when 3976 => b:="3976";
                when 3977 => b:="3977";
                when 3978 => b:="3978";
                when 3979 => b:="3979";
                when 3980 => b:="3980";
                when 3981 => b:="3981";
                when 3982 => b:="3982";
                when 3983 => b:="3983";
                when 3984 => b:="3984";
                when 3985 => b:="3985";
                when 3986 => b:="3986";
                when 3987 => b:="3987";
                when 3988 => b:="3988";
                when 3989 => b:="3989";
                when 3990 => b:="3990";
                when 3991 => b:="3991";
                when 3992 => b:="3992";
                when 3993 => b:="3993";
                when 3994 => b:="3994";
                when 3995 => b:="3995";
                when 3996 => b:="3996";
                when 3997 => b:="3997";
                when 3998 => b:="3998";
                when 4000 => b:="4000";
                when 4001 => b:="4001";
                when 4002 => b:="4002";
                when 4003 => b:="4003";
                when 4004 => b:="4004";
                when 4005 => b:="4005";
                when 4006 => b:="4006";
                when 4007 => b:="4007";
                when 4008 => b:="4008";
                when 4009 => b:="4009";
                when 4010 => b:="4010";
                when 4011 => b:="4011";
                when 4012 => b:="4012";
                when 4013 => b:="4013";
                when 4014 => b:="4014";
                when 4015 => b:="4015";
                when 4016 => b:="4016";
                when 4017 => b:="4017";
                when 4018 => b:="4018";
                when 4019 => b:="4019";
                when 4020 => b:="4020";
                when 4021 => b:="4021";
                when 4022 => b:="4022";
                when 4023 => b:="4023";
                when 4024 => b:="4024";
                when 4025 => b:="4025";
                when 4026 => b:="4026";
                when 4027 => b:="4027";
                when 4028 => b:="4028";
                when 4029 => b:="4029";
                when 4030 => b:="4030";
                when 4031 => b:="4031";
                when 4032 => b:="4032";
                when 4033 => b:="4033";
                when 4034 => b:="4034";
                when 4035 => b:="4035";
                when 4036 => b:="4036";
                when 4037 => b:="4037";
                when 4038 => b:="4038";
                when 4039 => b:="4039";
                when 4040 => b:="4040";
                when 4041 => b:="4041";
                when 4042 => b:="4042";
                when 4043 => b:="4043";
                when 4044 => b:="4044";
                when 4045 => b:="4045";
                when 4046 => b:="4046";
                when 4047 => b:="4047";
                when 4048 => b:="4048";
                when 4049 => b:="4049";
                when 4050 => b:="4050";
                when 4051 => b:="4051";
                when 4052 => b:="4052";
                when 4053 => b:="4053";
                when 4054 => b:="4054";
                when 4055 => b:="4055";
                when 4056 => b:="4056";
                when 4057 => b:="4057";
                when 4058 => b:="4058";
                when 4059 => b:="4059";
                when 4060 => b:="4060";
                when 4061 => b:="4061";
                when 4062 => b:="4062";
                when 4063 => b:="4063";
                when 4064 => b:="4064";
                when 4065 => b:="4065";
                when 4066 => b:="4066";
                when 4067 => b:="4067";
                when 4068 => b:="4068";
                when 4069 => b:="4069";
                when 4070 => b:="4070";
                when 4071 => b:="4071";
                when 4072 => b:="4072";
                when 4073 => b:="4073";
                when 4074 => b:="4074";
                when 4075 => b:="4075";
                when 4076 => b:="4076";
                when 4077 => b:="4077";
                when 4078 => b:="4078";
                when 4079 => b:="4079";
                when 4080 => b:="4080";
                when 4081 => b:="4081";
                when 4082 => b:="4082";
                when 4083 => b:="4083";
                when 4084 => b:="4084";
                when 4085 => b:="4085";
                when 4086 => b:="4086";
                when 4087 => b:="4087";
                when 4088 => b:="4088";
                when 4089 => b:="4089";
                when 4090 => b:="4090";
                when 4091 => b:="4091";
                when 4092 => b:="4092";
                when 4093 => b:="4093";
                when 4094 => b:="4094";
                when 4095 => b:="4095";
                when 4096 => b:="4096";
                when 4097 => b:="4097";
                when 4098 => b:="4098";
                when 4099 => b:="4099";
                when 4100 => b:="4100";
                when 4101 => b:="4101";
                when 4102 => b:="4102";
                when 4103 => b:="4103";
                when 4104 => b:="4104";
                when 4105 => b:="4105";
                when 4106 => b:="4106";
                when 4107 => b:="4107";
                when 4108 => b:="4108";
                when 4109 => b:="4109";
                when 4110 => b:="4110";
                when 4111 => b:="4111";
                when 4112 => b:="4112";
                when 4113 => b:="4113";
                when 4114 => b:="4114";
                when 4115 => b:="4115";
                when 4116 => b:="4116";
                when 4117 => b:="4117";
                when 4118 => b:="4118";
                when 4119 => b:="4119";
                when 4120 => b:="4120";
                when 4121 => b:="4121";
                when 4122 => b:="4122";
                when 4123 => b:="4123";
                when 4124 => b:="4124";
                when 4125 => b:="4125";
                when 4126 => b:="4126";
                when 4127 => b:="4127";
                when 4128 => b:="4128";
                when 4129 => b:="4129";
                when 4130 => b:="4130";
                when 4131 => b:="4131";
                when 4132 => b:="4132";
                when 4133 => b:="4133";
                when 4134 => b:="4134";
                when 4135 => b:="4135";
                when 4136 => b:="4136";
                when 4137 => b:="4137";
                when 4138 => b:="4138";
                when 4139 => b:="4139";
                when 4140 => b:="4140";
                when 4141 => b:="4141";
                when 4142 => b:="4142";
                when 4143 => b:="4143";
                when 4144 => b:="4144";
                when 4145 => b:="4145";
                when 4146 => b:="4146";
                when 4147 => b:="4147";
                when 4148 => b:="4148";
                when 4149 => b:="4149";
                when 4150 => b:="4150";
                when 4151 => b:="4151";
                when 4152 => b:="4152";
                when 4153 => b:="4153";
                when 4154 => b:="4154";
                when 4155 => b:="4155";
                when 4156 => b:="4156";
                when 4157 => b:="4157";
                when 4158 => b:="4158";
                when 4159 => b:="4159";
                when 4160 => b:="4160";
                when 4161 => b:="4161";
                when 4162 => b:="4162";
                when 4163 => b:="4163";
                when 4164 => b:="4164";
                when 4165 => b:="4165";
                when 4166 => b:="4166";
                when 4167 => b:="4167";
                when 4168 => b:="4168";
                when 4169 => b:="4169";
                when 4170 => b:="4170";
                when 4171 => b:="4171";
                when 4172 => b:="4172";
                when 4173 => b:="4173";
                when 4174 => b:="4174";
                when 4175 => b:="4175";
                when 4176 => b:="4176";
                when 4177 => b:="4177";
                when 4178 => b:="4178";
                when 4179 => b:="4179";
                when 4180 => b:="4180";
                when 4181 => b:="4181";
                when 4182 => b:="4182";
                when 4183 => b:="4183";
                when 4184 => b:="4184";
                when 4185 => b:="4185";
                when 4186 => b:="4186";
                when 4187 => b:="4187";
                when 4188 => b:="4188";
                when 4189 => b:="4189";
                when 4190 => b:="4190";
                when 4191 => b:="4191";
                when 4192 => b:="4192";
                when 4193 => b:="4193";
                when 4194 => b:="4194";
                when 4195 => b:="4195";
                when 4196 => b:="4196";
                when 4197 => b:="4197";
                when 4198 => b:="4198";
                when 4199 => b:="4199";
                when 4200 => b:="4200";
                when 4201 => b:="4201";
                when 4202 => b:="4202";
                when 4203 => b:="4203";
                when 4204 => b:="4204";
                when 4205 => b:="4205";
                when 4206 => b:="4206";
                when 4207 => b:="4207";
                when 4208 => b:="4208";
                when 4209 => b:="4209";
                when 4210 => b:="4210";
                when 4211 => b:="4211";
                when 4212 => b:="4212";
                when 4213 => b:="4213";
                when 4214 => b:="4214";
                when 4215 => b:="4215";
                when 4216 => b:="4216";
                when 4217 => b:="4217";
                when 4218 => b:="4218";
                when 4219 => b:="4219";
                when 4220 => b:="4220";
                when 4221 => b:="4221";
                when 4222 => b:="4222";
                when 4223 => b:="4223";
                when 4224 => b:="4224";
                when 4225 => b:="4225";
                when 4226 => b:="4226";
                when 4227 => b:="4227";
                when 4228 => b:="4228";
                when 4229 => b:="4229";
                when 4230 => b:="4230";
                when 4231 => b:="4231";
                when 4232 => b:="4232";
                when 4233 => b:="4233";
                when 4234 => b:="4234";
                when 4235 => b:="4235";
                when 4236 => b:="4236";
                when 4237 => b:="4237";
                when 4238 => b:="4238";
                when 4239 => b:="4239";
                when 4240 => b:="4240";
                when 4241 => b:="4241";
                when 4242 => b:="4242";
                when 4243 => b:="4243";
                when 4244 => b:="4244";
                when 4245 => b:="4245";
                when 4246 => b:="4246";
                when 4247 => b:="4247";
                when 4248 => b:="4248";
                when 4249 => b:="4249";
                when 4250 => b:="4250";
                when 4251 => b:="4251";
                when 4252 => b:="4252";
                when 4253 => b:="4253";
                when 4254 => b:="4254";
                when 4255 => b:="4255";
                when 4256 => b:="4256";
                when 4257 => b:="4257";
                when 4258 => b:="4258";
                when 4259 => b:="4259";
                when 4260 => b:="4260";
                when 4261 => b:="4261";
                when 4262 => b:="4262";
                when 4263 => b:="4263";
                when 4264 => b:="4264";
                when 4265 => b:="4265";
                when 4266 => b:="4266";
                when 4267 => b:="4267";
                when 4268 => b:="4268";
                when 4269 => b:="4269";
                when 4270 => b:="4270";
                when 4271 => b:="4271";
                when 4272 => b:="4272";
                when 4273 => b:="4273";
                when 4274 => b:="4274";
                when 4275 => b:="4275";
                when 4276 => b:="4276";
                when 4277 => b:="4277";
                when 4278 => b:="4278";
                when 4279 => b:="4279";
                when 4280 => b:="4280";
                when 4281 => b:="4281";
                when 4282 => b:="4282";
                when 4283 => b:="4283";
                when 4284 => b:="4284";
                when 4285 => b:="4285";
                when 4286 => b:="4286";
                when 4287 => b:="4287";
                when 4288 => b:="4288";
                when 4289 => b:="4289";
                when 4290 => b:="4290";
                when 4291 => b:="4291";
                when 4292 => b:="4292";
                when 4293 => b:="4293";
                when 4294 => b:="4294";
                when 4295 => b:="4295";
                when 4296 => b:="4296";
                when 4297 => b:="4297";
                when 4298 => b:="4298";
                when 4299 => b:="4299";
                when 4300 => b:="4300";
                when 4301 => b:="4301";
                when 4302 => b:="4302";
                when 4303 => b:="4303";
                when 4304 => b:="4304";
                when 4305 => b:="4305";
                when 4306 => b:="4306";
                when 4307 => b:="4307";
                when 4308 => b:="4308";
                when 4309 => b:="4309";
                when 4310 => b:="4310";
                when 4311 => b:="4311";
                when 4312 => b:="4312";
                when 4313 => b:="4313";
                when 4314 => b:="4314";
                when 4315 => b:="4315";
                when 4316 => b:="4316";
                when 4317 => b:="4317";
                when 4318 => b:="4318";
                when 4319 => b:="4319";
                when 4320 => b:="4320";
                when 4321 => b:="4321";
                when 4322 => b:="4322";
                when 4323 => b:="4323";
                when 4324 => b:="4324";
                when 4325 => b:="4325";
                when 4326 => b:="4326";
                when 4327 => b:="4327";
                when 4328 => b:="4328";
                when 4329 => b:="4329";
                when 4330 => b:="4330";
                when 4331 => b:="4331";
                when 4332 => b:="4332";
                when 4333 => b:="4333";
                when 4334 => b:="4334";
                when 4335 => b:="4335";
                when 4336 => b:="4336";
                when 4337 => b:="4337";
                when 4338 => b:="4338";
                when 4339 => b:="4339";
                when 4340 => b:="4340";
                when 4341 => b:="4341";
                when 4342 => b:="4342";
                when 4343 => b:="4343";
                when 4344 => b:="4344";
                when 4345 => b:="4345";
                when 4346 => b:="4346";
                when 4347 => b:="4347";
                when 4348 => b:="4348";
                when 4349 => b:="4349";
                when 4350 => b:="4350";
                when 4351 => b:="4351";
                when 4352 => b:="4352";
                when 4353 => b:="4353";
                when 4354 => b:="4354";
                when 4355 => b:="4355";
                when 4356 => b:="4356";
                when 4357 => b:="4357";
                when 4358 => b:="4358";
                when 4359 => b:="4359";
                when 4360 => b:="4360";
                when 4361 => b:="4361";
                when 4362 => b:="4362";
                when 4363 => b:="4363";
                when 4364 => b:="4364";
                when 4365 => b:="4365";
                when 4366 => b:="4366";
                when 4367 => b:="4367";
                when 4368 => b:="4368";
                when 4369 => b:="4369";
                when 4370 => b:="4370";
                when 4371 => b:="4371";
                when 4372 => b:="4372";
                when 4373 => b:="4373";
                when 4374 => b:="4374";
                when 4375 => b:="4375";
                when 4376 => b:="4376";
                when 4377 => b:="4377";
                when 4378 => b:="4378";
                when 4379 => b:="4379";
                when 4380 => b:="4380";
                when 4381 => b:="4381";
                when 4382 => b:="4382";
                when 4383 => b:="4383";
                when 4384 => b:="4384";
                when 4385 => b:="4385";
                when 4386 => b:="4386";
                when 4387 => b:="4387";
                when 4388 => b:="4388";
                when 4389 => b:="4389";
                when 4390 => b:="4390";
                when 4391 => b:="4391";
                when 4392 => b:="4392";
                when 4393 => b:="4393";
                when 4394 => b:="4394";
                when 4395 => b:="4395";
                when 4396 => b:="4396";
                when 4397 => b:="4397";
                when 4398 => b:="4398";
                when 4399 => b:="4399";
                when 4400 => b:="4400";
                when 4401 => b:="4401";
                when 4402 => b:="4402";
                when 4403 => b:="4403";
                when 4404 => b:="4404";
                when 4405 => b:="4405";
                when 4406 => b:="4406";
                when 4407 => b:="4407";
                when 4408 => b:="4408";
                when 4409 => b:="4409";
                when 4410 => b:="4410";
                when 4411 => b:="4411";
                when 4412 => b:="4412";
                when 4413 => b:="4413";
                when 4414 => b:="4414";
                when 4415 => b:="4415";
                when 4416 => b:="4416";
                when 4417 => b:="4417";
                when 4418 => b:="4418";
                when 4419 => b:="4419";
                when 4420 => b:="4420";
                when 4421 => b:="4421";
                when 4422 => b:="4422";
                when 4423 => b:="4423";
                when 4424 => b:="4424";
                when 4425 => b:="4425";
                when 4426 => b:="4426";
                when 4427 => b:="4427";
                when 4428 => b:="4428";
                when 4429 => b:="4429";
                when 4430 => b:="4430";
                when 4431 => b:="4431";
                when 4432 => b:="4432";
                when 4433 => b:="4433";
                when 4434 => b:="4434";
                when 4435 => b:="4435";
                when 4436 => b:="4436";
                when 4437 => b:="4437";
                when 4438 => b:="4438";
                when 4439 => b:="4439";
                when 4440 => b:="4440";
                when 4441 => b:="4441";
                when 4442 => b:="4442";
                when 4443 => b:="4443";
                when 4444 => b:="4444";
                when 4445 => b:="4445";
                when 4446 => b:="4446";
                when 4447 => b:="4447";
                when 4448 => b:="4448";
                when 4449 => b:="4449";
                when 4450 => b:="4450";
                when 4451 => b:="4451";
                when 4452 => b:="4452";
                when 4453 => b:="4453";
                when 4454 => b:="4454";
                when 4455 => b:="4455";
                when 4456 => b:="4456";
                when 4457 => b:="4457";
                when 4458 => b:="4458";
                when 4459 => b:="4459";
                when 4460 => b:="4460";
                when 4461 => b:="4461";
                when 4462 => b:="4462";
                when 4463 => b:="4463";
                when 4464 => b:="4464";
                when 4465 => b:="4465";
                when 4466 => b:="4466";
                when 4467 => b:="4467";
                when 4468 => b:="4468";
                when 4469 => b:="4469";
                when 4470 => b:="4470";
                when 4471 => b:="4471";
                when 4472 => b:="4472";
                when 4473 => b:="4473";
                when 4474 => b:="4474";
                when 4475 => b:="4475";
                when 4476 => b:="4476";
                when 4477 => b:="4477";
                when 4478 => b:="4478";
                when 4479 => b:="4479";
                when 4480 => b:="4480";
                when 4481 => b:="4481";
                when 4482 => b:="4482";
                when 4483 => b:="4483";
                when 4484 => b:="4484";
                when 4485 => b:="4485";
                when 4486 => b:="4486";
                when 4487 => b:="4487";
                when 4488 => b:="4488";
                when 4489 => b:="4489";
                when 4490 => b:="4490";
                when 4491 => b:="4491";
                when 4492 => b:="4492";
                when 4493 => b:="4493";
                when 4494 => b:="4494";
                when 4495 => b:="4495";
                when 4496 => b:="4496";
                when 4497 => b:="4497";
                when 4498 => b:="4498";
                when 4499 => b:="4499";
                when 4500 => b:="4500";
                when 4501 => b:="4501";
                when 4502 => b:="4502";
                when 4503 => b:="4503";
                when 4504 => b:="4504";
                when 4505 => b:="4505";
                when 4506 => b:="4506";
                when 4507 => b:="4507";
                when 4508 => b:="4508";
                when 4509 => b:="4509";
                when 4510 => b:="4510";
                when 4511 => b:="4511";
                when 4512 => b:="4512";
                when 4513 => b:="4513";
                when 4514 => b:="4514";
                when 4515 => b:="4515";
                when 4516 => b:="4516";
                when 4517 => b:="4517";
                when 4518 => b:="4518";
                when 4519 => b:="4519";
                when 4520 => b:="4520";
                when 4521 => b:="4521";
                when 4522 => b:="4522";
                when 4523 => b:="4523";
                when 4524 => b:="4524";
                when 4525 => b:="4525";
                when 4526 => b:="4526";
                when 4527 => b:="4527";
                when 4528 => b:="4528";
                when 4529 => b:="4529";
                when 4530 => b:="4530";
                when 4531 => b:="4531";
                when 4532 => b:="4532";
                when 4533 => b:="4533";
                when 4534 => b:="4534";
                when 4535 => b:="4535";
                when 4536 => b:="4536";
                when 4537 => b:="4537";
                when 4538 => b:="4538";
                when 4539 => b:="4539";
                when 4540 => b:="4540";
                when 4541 => b:="4541";
                when 4542 => b:="4542";
                when 4543 => b:="4543";
                when 4544 => b:="4544";
                when 4545 => b:="4545";
                when 4546 => b:="4546";
                when 4547 => b:="4547";
                when 4548 => b:="4548";
                when 4549 => b:="4549";
                when 4550 => b:="4550";
                when 4551 => b:="4551";
                when 4552 => b:="4552";
                when 4553 => b:="4553";
                when 4554 => b:="4554";
                when 4555 => b:="4555";
                when 4556 => b:="4556";
                when 4557 => b:="4557";
                when 4558 => b:="4558";
                when 4559 => b:="4559";
                when 4560 => b:="4560";
                when 4561 => b:="4561";
                when 4562 => b:="4562";
                when 4563 => b:="4563";
                when 4564 => b:="4564";
                when 4565 => b:="4565";
                when 4566 => b:="4566";
                when 4567 => b:="4567";
                when 4568 => b:="4568";
                when 4569 => b:="4569";
                when 4570 => b:="4570";
                when 4571 => b:="4571";
                when 4572 => b:="4572";
                when 4573 => b:="4573";
                when 4574 => b:="4574";
                when 4575 => b:="4575";
                when 4576 => b:="4576";
                when 4577 => b:="4577";
                when 4578 => b:="4578";
                when 4579 => b:="4579";
                when 4580 => b:="4580";
                when 4581 => b:="4581";
                when 4582 => b:="4582";
                when 4583 => b:="4583";
                when 4584 => b:="4584";
                when 4585 => b:="4585";
                when 4586 => b:="4586";
                when 4587 => b:="4587";
                when 4588 => b:="4588";
                when 4589 => b:="4589";
                when 4590 => b:="4590";
                when 4591 => b:="4591";
                when 4592 => b:="4592";
                when 4593 => b:="4593";
                when 4594 => b:="4594";
                when 4595 => b:="4595";
                when 4596 => b:="4596";
                when 4597 => b:="4597";
                when 4598 => b:="4598";
                when 4599 => b:="4599";
                when 4600 => b:="4600";
                when 4601 => b:="4601";
                when 4602 => b:="4602";
                when 4603 => b:="4603";
                when 4604 => b:="4604";
                when 4605 => b:="4605";
                when 4606 => b:="4606";
                when 4607 => b:="4607";
                when 4608 => b:="4608";
                when 4609 => b:="4609";
                when 4610 => b:="4610";
                when 4611 => b:="4611";
                when 4612 => b:="4612";
                when 4613 => b:="4613";
                when 4614 => b:="4614";
                when 4615 => b:="4615";
                when 4616 => b:="4616";
                when 4617 => b:="4617";
                when 4618 => b:="4618";
                when 4619 => b:="4619";
                when 4620 => b:="4620";
                when 4621 => b:="4621";
                when 4622 => b:="4622";
                when 4623 => b:="4623";
                when 4624 => b:="4624";
                when 4625 => b:="4625";
                when 4626 => b:="4626";
                when 4627 => b:="4627";
                when 4628 => b:="4628";
                when 4629 => b:="4629";
                when 4630 => b:="4630";
                when 4631 => b:="4631";
                when 4632 => b:="4632";
                when 4633 => b:="4633";
                when 4634 => b:="4634";
                when 4635 => b:="4635";
                when 4636 => b:="4636";
                when 4637 => b:="4637";
                when 4638 => b:="4638";
                when 4639 => b:="4639";
                when 4640 => b:="4640";
                when 4641 => b:="4641";
                when 4642 => b:="4642";
                when 4643 => b:="4643";
                when 4644 => b:="4644";
                when 4645 => b:="4645";
                when 4646 => b:="4646";
                when 4647 => b:="4647";
                when 4648 => b:="4648";
                when 4649 => b:="4649";
                when 4650 => b:="4650";
                when 4651 => b:="4651";
                when 4652 => b:="4652";
                when 4653 => b:="4653";
                when 4654 => b:="4654";
                when 4655 => b:="4655";
                when 4656 => b:="4656";
                when 4657 => b:="4657";
                when 4658 => b:="4658";
                when 4659 => b:="4659";
                when 4660 => b:="4660";
                when 4661 => b:="4661";
                when 4662 => b:="4662";
                when 4663 => b:="4663";
                when 4664 => b:="4664";
                when 4665 => b:="4665";
                when 4666 => b:="4666";
                when 4667 => b:="4667";
                when 4668 => b:="4668";
                when 4669 => b:="4669";
                when 4670 => b:="4670";
                when 4671 => b:="4671";
                when 4672 => b:="4672";
                when 4673 => b:="4673";
                when 4674 => b:="4674";
                when 4675 => b:="4675";
                when 4676 => b:="4676";
                when 4677 => b:="4677";
                when 4678 => b:="4678";
                when 4679 => b:="4679";
                when 4680 => b:="4680";
                when 4681 => b:="4681";
                when 4682 => b:="4682";
                when 4683 => b:="4683";
                when 4684 => b:="4684";
                when 4685 => b:="4685";
                when 4686 => b:="4686";
                when 4687 => b:="4687";
                when 4688 => b:="4688";
                when 4689 => b:="4689";
                when 4690 => b:="4690";
                when 4691 => b:="4691";
                when 4692 => b:="4692";
                when 4693 => b:="4693";
                when 4694 => b:="4694";
                when 4695 => b:="4695";
                when 4696 => b:="4696";
                when 4697 => b:="4697";
                when 4698 => b:="4698";
                when 4699 => b:="4699";
                when 4700 => b:="4700";
                when 4701 => b:="4701";
                when 4702 => b:="4702";
                when 4703 => b:="4703";
                when 4704 => b:="4704";
                when 4705 => b:="4705";
                when 4706 => b:="4706";
                when 4707 => b:="4707";
                when 4708 => b:="4708";
                when 4709 => b:="4709";
                when 4710 => b:="4710";
                when 4711 => b:="4711";
                when 4712 => b:="4712";
                when 4713 => b:="4713";
                when 4714 => b:="4714";
                when 4715 => b:="4715";
                when 4716 => b:="4716";
                when 4717 => b:="4717";
                when 4718 => b:="4718";
                when 4719 => b:="4719";
                when 4720 => b:="4720";
                when 4721 => b:="4721";
                when 4722 => b:="4722";
                when 4723 => b:="4723";
                when 4724 => b:="4724";
                when 4725 => b:="4725";
                when 4726 => b:="4726";
                when 4727 => b:="4727";
                when 4728 => b:="4728";
                when 4729 => b:="4729";
                when 4730 => b:="4730";
                when 4731 => b:="4731";
                when 4732 => b:="4732";
                when 4733 => b:="4733";
                when 4734 => b:="4734";
                when 4735 => b:="4735";
                when 4736 => b:="4736";
                when 4737 => b:="4737";
                when 4738 => b:="4738";
                when 4739 => b:="4739";
                when 4740 => b:="4740";
                when 4741 => b:="4741";
                when 4742 => b:="4742";
                when 4743 => b:="4743";
                when 4744 => b:="4744";
                when 4745 => b:="4745";
                when 4746 => b:="4746";
                when 4747 => b:="4747";
                when 4748 => b:="4748";
                when 4749 => b:="4749";
                when 4750 => b:="4750";
                when 4751 => b:="4751";
                when 4752 => b:="4752";
                when 4753 => b:="4753";
                when 4754 => b:="4754";
                when 4755 => b:="4755";
                when 4756 => b:="4756";
                when 4757 => b:="4757";
                when 4758 => b:="4758";
                when 4759 => b:="4759";
                when 4760 => b:="4760";
                when 4761 => b:="4761";
                when 4762 => b:="4762";
                when 4763 => b:="4763";
                when 4764 => b:="4764";
                when 4765 => b:="4765";
                when 4766 => b:="4766";
                when 4767 => b:="4767";
                when 4768 => b:="4768";
                when 4769 => b:="4769";
                when 4770 => b:="4770";
                when 4771 => b:="4771";
                when 4772 => b:="4772";
                when 4773 => b:="4773";
                when 4774 => b:="4774";
                when 4775 => b:="4775";
                when 4776 => b:="4776";
                when 4777 => b:="4777";
                when 4778 => b:="4778";
                when 4779 => b:="4779";
                when 4780 => b:="4780";
                when 4781 => b:="4781";
                when 4782 => b:="4782";
                when 4783 => b:="4783";
                when 4784 => b:="4784";
                when 4785 => b:="4785";
                when 4786 => b:="4786";
                when 4787 => b:="4787";
                when 4788 => b:="4788";
                when 4789 => b:="4789";
                when 4790 => b:="4790";
                when 4791 => b:="4791";
                when 4792 => b:="4792";
                when 4793 => b:="4793";
                when 4794 => b:="4794";
                when 4795 => b:="4795";
                when 4796 => b:="4796";
                when 4797 => b:="4797";
                when 4798 => b:="4798";
                when 4799 => b:="4799";
                when 4800 => b:="4800";
                when 4801 => b:="4801";
                when 4802 => b:="4802";
                when 4803 => b:="4803";
                when 4804 => b:="4804";
                when 4805 => b:="4805";
                when 4806 => b:="4806";
                when 4807 => b:="4807";
                when 4808 => b:="4808";
                when 4809 => b:="4809";
                when 4810 => b:="4810";
                when 4811 => b:="4811";
                when 4812 => b:="4812";
                when 4813 => b:="4813";
                when 4814 => b:="4814";
                when 4815 => b:="4815";
                when 4816 => b:="4816";
                when 4817 => b:="4817";
                when 4818 => b:="4818";
                when 4819 => b:="4819";
                when 4820 => b:="4820";
                when 4821 => b:="4821";
                when 4822 => b:="4822";
                when 4823 => b:="4823";
                when 4824 => b:="4824";
                when 4825 => b:="4825";
                when 4826 => b:="4826";
                when 4827 => b:="4827";
                when 4828 => b:="4828";
                when 4829 => b:="4829";
                when 4830 => b:="4830";
                when 4831 => b:="4831";
                when 4832 => b:="4832";
                when 4833 => b:="4833";
                when 4834 => b:="4834";
                when 4835 => b:="4835";
                when 4836 => b:="4836";
                when 4837 => b:="4837";
                when 4838 => b:="4838";
                when 4839 => b:="4839";
                when 4840 => b:="4840";
                when 4841 => b:="4841";
                when 4842 => b:="4842";
                when 4843 => b:="4843";
                when 4844 => b:="4844";
                when 4845 => b:="4845";
                when 4846 => b:="4846";
                when 4847 => b:="4847";
                when 4848 => b:="4848";
                when 4849 => b:="4849";
                when 4850 => b:="4850";
                when 4851 => b:="4851";
                when 4852 => b:="4852";
                when 4853 => b:="4853";
                when 4854 => b:="4854";
                when 4855 => b:="4855";
                when 4856 => b:="4856";
                when 4857 => b:="4857";
                when 4858 => b:="4858";
                when 4859 => b:="4859";
                when 4860 => b:="4860";
                when 4861 => b:="4861";
                when 4862 => b:="4862";
                when 4863 => b:="4863";
                when 4864 => b:="4864";
                when 4865 => b:="4865";
                when 4866 => b:="4866";
                when 4867 => b:="4867";
                when 4868 => b:="4868";
                when 4869 => b:="4869";
                when 4870 => b:="4870";
                when 4871 => b:="4871";
                when 4872 => b:="4872";
                when 4873 => b:="4873";
                when 4874 => b:="4874";
                when 4875 => b:="4875";
                when 4876 => b:="4876";
                when 4877 => b:="4877";
                when 4878 => b:="4878";
                when 4879 => b:="4879";
                when 4880 => b:="4880";
                when 4881 => b:="4881";
                when 4882 => b:="4882";
                when 4883 => b:="4883";
                when 4884 => b:="4884";
                when 4885 => b:="4885";
                when 4886 => b:="4886";
                when 4887 => b:="4887";
                when 4888 => b:="4888";
                when 4889 => b:="4889";
                when 4890 => b:="4890";
                when 4891 => b:="4891";
                when 4892 => b:="4892";
                when 4893 => b:="4893";
                when 4894 => b:="4894";
                when 4895 => b:="4895";
                when 4896 => b:="4896";
                when 4897 => b:="4897";
                when 4898 => b:="4898";
                when 4899 => b:="4899";
                when 4900 => b:="4900";
                when 4901 => b:="4901";
                when 4902 => b:="4902";
                when 4903 => b:="4903";
                when 4904 => b:="4904";
                when 4905 => b:="4905";
                when 4906 => b:="4906";
                when 4907 => b:="4907";
                when 4908 => b:="4908";
                when 4909 => b:="4909";
                when 4910 => b:="4910";
                when 4911 => b:="4911";
                when 4912 => b:="4912";
                when 4913 => b:="4913";
                when 4914 => b:="4914";
                when 4915 => b:="4915";
                when 4916 => b:="4916";
                when 4917 => b:="4917";
                when 4918 => b:="4918";
                when 4919 => b:="4919";
                when 4920 => b:="4920";
                when 4921 => b:="4921";
                when 4922 => b:="4922";
                when 4923 => b:="4923";
                when 4924 => b:="4924";
                when 4925 => b:="4925";
                when 4926 => b:="4926";
                when 4927 => b:="4927";
                when 4928 => b:="4928";
                when 4929 => b:="4929";
                when 4930 => b:="4930";
                when 4931 => b:="4931";
                when 4932 => b:="4932";
                when 4933 => b:="4933";
                when 4934 => b:="4934";
                when 4935 => b:="4935";
                when 4936 => b:="4936";
                when 4937 => b:="4937";
                when 4938 => b:="4938";
                when 4939 => b:="4939";
                when 4940 => b:="4940";
                when 4941 => b:="4941";
                when 4942 => b:="4942";
                when 4943 => b:="4943";
                when 4944 => b:="4944";
                when 4945 => b:="4945";
                when 4946 => b:="4946";
                when 4947 => b:="4947";
                when 4948 => b:="4948";
                when 4949 => b:="4949";
                when 4950 => b:="4950";
                when 4951 => b:="4951";
                when 4952 => b:="4952";
                when 4953 => b:="4953";
                when 4954 => b:="4954";
                when 4955 => b:="4955";
                when 4956 => b:="4956";
                when 4957 => b:="4957";
                when 4958 => b:="4958";
                when 4959 => b:="4959";
                when 4960 => b:="4960";
                when 4961 => b:="4961";
                when 4962 => b:="4962";
                when 4963 => b:="4963";
                when 4964 => b:="4964";
                when 4965 => b:="4965";
                when 4966 => b:="4966";
                when 4967 => b:="4967";
                when 4968 => b:="4968";
                when 4969 => b:="4969";
                when 4970 => b:="4970";
                when 4971 => b:="4971";
                when 4972 => b:="4972";
                when 4973 => b:="4973";
                when 4974 => b:="4974";
                when 4975 => b:="4975";
                when 4976 => b:="4976";
                when 4977 => b:="4977";
                when 4978 => b:="4978";
                when 4979 => b:="4979";
                when 4980 => b:="4980";
                when 4981 => b:="4981";
                when 4982 => b:="4982";
                when 4983 => b:="4983";
                when 4984 => b:="4984";
                when 4985 => b:="4985";
                when 4986 => b:="4986";
                when 4987 => b:="4987";
                when 4988 => b:="4988";
                when 4989 => b:="4989";
                when 4990 => b:="4990";
                when 4991 => b:="4991";
                when 4992 => b:="4992";
                when 4993 => b:="4993";
                when 4994 => b:="4994";
                when 4995 => b:="4995";
                when 4996 => b:="4996";
                when 4997 => b:="4997";
                when 4998 => b:="4998";
                when 5000 => b:="5000";
                when 5001 => b:="5001";
                when 5002 => b:="5002";
                when 5003 => b:="5003";
                when 5004 => b:="5004";
                when 5005 => b:="5005";
                when 5006 => b:="5006";
                when 5007 => b:="5007";
                when 5008 => b:="5008";
                when 5009 => b:="5009";
                when 5010 => b:="5010";
                when 5011 => b:="5011";
                when 5012 => b:="5012";
                when 5013 => b:="5013";
                when 5014 => b:="5014";
                when 5015 => b:="5015";
                when 5016 => b:="5016";
                when 5017 => b:="5017";
                when 5018 => b:="5018";
                when 5019 => b:="5019";
                when 5020 => b:="5020";
                when 5021 => b:="5021";
                when 5022 => b:="5022";
                when 5023 => b:="5023";
                when 5024 => b:="5024";
                when 5025 => b:="5025";
                when 5026 => b:="5026";
                when 5027 => b:="5027";
                when 5028 => b:="5028";
                when 5029 => b:="5029";
                when 5030 => b:="5030";
                when 5031 => b:="5031";
                when 5032 => b:="5032";
                when 5033 => b:="5033";
                when 5034 => b:="5034";
                when 5035 => b:="5035";
                when 5036 => b:="5036";
                when 5037 => b:="5037";
                when 5038 => b:="5038";
                when 5039 => b:="5039";
                when 5040 => b:="5040";
                when 5041 => b:="5041";
                when 5042 => b:="5042";
                when 5043 => b:="5043";
                when 5044 => b:="5044";
                when 5045 => b:="5045";
                when 5046 => b:="5046";
                when 5047 => b:="5047";
                when 5048 => b:="5048";
                when 5049 => b:="5049";
                when 5050 => b:="5050";
                when 5051 => b:="5051";
                when 5052 => b:="5052";
                when 5053 => b:="5053";
                when 5054 => b:="5054";
                when 5055 => b:="5055";
                when 5056 => b:="5056";
                when 5057 => b:="5057";
                when 5058 => b:="5058";
                when 5059 => b:="5059";
                when 5060 => b:="5060";
                when 5061 => b:="5061";
                when 5062 => b:="5062";
                when 5063 => b:="5063";
                when 5064 => b:="5064";
                when 5065 => b:="5065";
                when 5066 => b:="5066";
                when 5067 => b:="5067";
                when 5068 => b:="5068";
                when 5069 => b:="5069";
                when 5070 => b:="5070";
                when 5071 => b:="5071";
                when 5072 => b:="5072";
                when 5073 => b:="5073";
                when 5074 => b:="5074";
                when 5075 => b:="5075";
                when 5076 => b:="5076";
                when 5077 => b:="5077";
                when 5078 => b:="5078";
                when 5079 => b:="5079";
                when 5080 => b:="5080";
                when 5081 => b:="5081";
                when 5082 => b:="5082";
                when 5083 => b:="5083";
                when 5084 => b:="5084";
                when 5085 => b:="5085";
                when 5086 => b:="5086";
                when 5087 => b:="5087";
                when 5088 => b:="5088";
                when 5089 => b:="5089";
                when 5090 => b:="5090";
                when 5091 => b:="5091";
                when 5092 => b:="5092";
                when 5093 => b:="5093";
                when 5094 => b:="5094";
                when 5095 => b:="5095";
                when 5096 => b:="5096";
                when 5097 => b:="5097";
                when 5098 => b:="5098";
                when 5099 => b:="5099";
                when 5100 => b:="5100";
                when 5101 => b:="5101";
                when 5102 => b:="5102";
                when 5103 => b:="5103";
                when 5104 => b:="5104";
                when 5105 => b:="5105";
                when 5106 => b:="5106";
                when 5107 => b:="5107";
                when 5108 => b:="5108";
                when 5109 => b:="5109";
                when 5110 => b:="5110";
                when 5111 => b:="5111";
                when 5112 => b:="5112";
                when 5113 => b:="5113";
                when 5114 => b:="5114";
                when 5115 => b:="5115";
                when 5116 => b:="5116";
                when 5117 => b:="5117";
                when 5118 => b:="5118";
                when 5119 => b:="5119";
                when 5120 => b:="5120";
                when 5121 => b:="5121";
                when 5122 => b:="5122";
                when 5123 => b:="5123";
                when 5124 => b:="5124";
                when 5125 => b:="5125";
                when 5126 => b:="5126";
                when 5127 => b:="5127";
                when 5128 => b:="5128";
                when 5129 => b:="5129";
                when 5130 => b:="5130";
                when 5131 => b:="5131";
                when 5132 => b:="5132";
                when 5133 => b:="5133";
                when 5134 => b:="5134";
                when 5135 => b:="5135";
                when 5136 => b:="5136";
                when 5137 => b:="5137";
                when 5138 => b:="5138";
                when 5139 => b:="5139";
                when 5140 => b:="5140";
                when 5141 => b:="5141";
                when 5142 => b:="5142";
                when 5143 => b:="5143";
                when 5144 => b:="5144";
                when 5145 => b:="5145";
                when 5146 => b:="5146";
                when 5147 => b:="5147";
                when 5148 => b:="5148";
                when 5149 => b:="5149";
                when 5150 => b:="5150";
                when 5151 => b:="5151";
                when 5152 => b:="5152";
                when 5153 => b:="5153";
                when 5154 => b:="5154";
                when 5155 => b:="5155";
                when 5156 => b:="5156";
                when 5157 => b:="5157";
                when 5158 => b:="5158";
                when 5159 => b:="5159";
                when 5160 => b:="5160";
                when 5161 => b:="5161";
                when 5162 => b:="5162";
                when 5163 => b:="5163";
                when 5164 => b:="5164";
                when 5165 => b:="5165";
                when 5166 => b:="5166";
                when 5167 => b:="5167";
                when 5168 => b:="5168";
                when 5169 => b:="5169";
                when 5170 => b:="5170";
                when 5171 => b:="5171";
                when 5172 => b:="5172";
                when 5173 => b:="5173";
                when 5174 => b:="5174";
                when 5175 => b:="5175";
                when 5176 => b:="5176";
                when 5177 => b:="5177";
                when 5178 => b:="5178";
                when 5179 => b:="5179";
                when 5180 => b:="5180";
                when 5181 => b:="5181";
                when 5182 => b:="5182";
                when 5183 => b:="5183";
                when 5184 => b:="5184";
                when 5185 => b:="5185";
                when 5186 => b:="5186";
                when 5187 => b:="5187";
                when 5188 => b:="5188";
                when 5189 => b:="5189";
                when 5190 => b:="5190";
                when 5191 => b:="5191";
                when 5192 => b:="5192";
                when 5193 => b:="5193";
                when 5194 => b:="5194";
                when 5195 => b:="5195";
                when 5196 => b:="5196";
                when 5197 => b:="5197";
                when 5198 => b:="5198";
                when 5199 => b:="5199";
                when 5200 => b:="5200";
                when 5201 => b:="5201";
                when 5202 => b:="5202";
                when 5203 => b:="5203";
                when 5204 => b:="5204";
                when 5205 => b:="5205";
                when 5206 => b:="5206";
                when 5207 => b:="5207";
                when 5208 => b:="5208";
                when 5209 => b:="5209";
                when 5210 => b:="5210";
                when 5211 => b:="5211";
                when 5212 => b:="5212";
                when 5213 => b:="5213";
                when 5214 => b:="5214";
                when 5215 => b:="5215";
                when 5216 => b:="5216";
                when 5217 => b:="5217";
                when 5218 => b:="5218";
                when 5219 => b:="5219";
                when 5220 => b:="5220";
                when 5221 => b:="5221";
                when 5222 => b:="5222";
                when 5223 => b:="5223";
                when 5224 => b:="5224";
                when 5225 => b:="5225";
                when 5226 => b:="5226";
                when 5227 => b:="5227";
                when 5228 => b:="5228";
                when 5229 => b:="5229";
                when 5230 => b:="5230";
                when 5231 => b:="5231";
                when 5232 => b:="5232";
                when 5233 => b:="5233";
                when 5234 => b:="5234";
                when 5235 => b:="5235";
                when 5236 => b:="5236";
                when 5237 => b:="5237";
                when 5238 => b:="5238";
                when 5239 => b:="5239";
                when 5240 => b:="5240";
                when 5241 => b:="5241";
                when 5242 => b:="5242";
                when 5243 => b:="5243";
                when 5244 => b:="5244";
                when 5245 => b:="5245";
                when 5246 => b:="5246";
                when 5247 => b:="5247";
                when 5248 => b:="5248";
                when 5249 => b:="5249";
                when 5250 => b:="5250";
                when 5251 => b:="5251";
                when 5252 => b:="5252";
                when 5253 => b:="5253";
                when 5254 => b:="5254";
                when 5255 => b:="5255";
                when 5256 => b:="5256";
                when 5257 => b:="5257";
                when 5258 => b:="5258";
                when 5259 => b:="5259";
                when 5260 => b:="5260";
                when 5261 => b:="5261";
                when 5262 => b:="5262";
                when 5263 => b:="5263";
                when 5264 => b:="5264";
                when 5265 => b:="5265";
                when 5266 => b:="5266";
                when 5267 => b:="5267";
                when 5268 => b:="5268";
                when 5269 => b:="5269";
                when 5270 => b:="5270";
                when 5271 => b:="5271";
                when 5272 => b:="5272";
                when 5273 => b:="5273";
                when 5274 => b:="5274";
                when 5275 => b:="5275";
                when 5276 => b:="5276";
                when 5277 => b:="5277";
                when 5278 => b:="5278";
                when 5279 => b:="5279";
                when 5280 => b:="5280";
                when 5281 => b:="5281";
                when 5282 => b:="5282";
                when 5283 => b:="5283";
                when 5284 => b:="5284";
                when 5285 => b:="5285";
                when 5286 => b:="5286";
                when 5287 => b:="5287";
                when 5288 => b:="5288";
                when 5289 => b:="5289";
                when 5290 => b:="5290";
                when 5291 => b:="5291";
                when 5292 => b:="5292";
                when 5293 => b:="5293";
                when 5294 => b:="5294";
                when 5295 => b:="5295";
                when 5296 => b:="5296";
                when 5297 => b:="5297";
                when 5298 => b:="5298";
                when 5299 => b:="5299";
                when 5300 => b:="5300";
                when 5301 => b:="5301";
                when 5302 => b:="5302";
                when 5303 => b:="5303";
                when 5304 => b:="5304";
                when 5305 => b:="5305";
                when 5306 => b:="5306";
                when 5307 => b:="5307";
                when 5308 => b:="5308";
                when 5309 => b:="5309";
                when 5310 => b:="5310";
                when 5311 => b:="5311";
                when 5312 => b:="5312";
                when 5313 => b:="5313";
                when 5314 => b:="5314";
                when 5315 => b:="5315";
                when 5316 => b:="5316";
                when 5317 => b:="5317";
                when 5318 => b:="5318";
                when 5319 => b:="5319";
                when 5320 => b:="5320";
                when 5321 => b:="5321";
                when 5322 => b:="5322";
                when 5323 => b:="5323";
                when 5324 => b:="5324";
                when 5325 => b:="5325";
                when 5326 => b:="5326";
                when 5327 => b:="5327";
                when 5328 => b:="5328";
                when 5329 => b:="5329";
                when 5330 => b:="5330";
                when 5331 => b:="5331";
                when 5332 => b:="5332";
                when 5333 => b:="5333";
                when 5334 => b:="5334";
                when 5335 => b:="5335";
                when 5336 => b:="5336";
                when 5337 => b:="5337";
                when 5338 => b:="5338";
                when 5339 => b:="5339";
                when 5340 => b:="5340";
                when 5341 => b:="5341";
                when 5342 => b:="5342";
                when 5343 => b:="5343";
                when 5344 => b:="5344";
                when 5345 => b:="5345";
                when 5346 => b:="5346";
                when 5347 => b:="5347";
                when 5348 => b:="5348";
                when 5349 => b:="5349";
                when 5350 => b:="5350";
                when 5351 => b:="5351";
                when 5352 => b:="5352";
                when 5353 => b:="5353";
                when 5354 => b:="5354";
                when 5355 => b:="5355";
                when 5356 => b:="5356";
                when 5357 => b:="5357";
                when 5358 => b:="5358";
                when 5359 => b:="5359";
                when 5360 => b:="5360";
                when 5361 => b:="5361";
                when 5362 => b:="5362";
                when 5363 => b:="5363";
                when 5364 => b:="5364";
                when 5365 => b:="5365";
                when 5366 => b:="5366";
                when 5367 => b:="5367";
                when 5368 => b:="5368";
                when 5369 => b:="5369";
                when 5370 => b:="5370";
                when 5371 => b:="5371";
                when 5372 => b:="5372";
                when 5373 => b:="5373";
                when 5374 => b:="5374";
                when 5375 => b:="5375";
                when 5376 => b:="5376";
                when 5377 => b:="5377";
                when 5378 => b:="5378";
                when 5379 => b:="5379";
                when 5380 => b:="5380";
                when 5381 => b:="5381";
                when 5382 => b:="5382";
                when 5383 => b:="5383";
                when 5384 => b:="5384";
                when 5385 => b:="5385";
                when 5386 => b:="5386";
                when 5387 => b:="5387";
                when 5388 => b:="5388";
                when 5389 => b:="5389";
                when 5390 => b:="5390";
                when 5391 => b:="5391";
                when 5392 => b:="5392";
                when 5393 => b:="5393";
                when 5394 => b:="5394";
                when 5395 => b:="5395";
                when 5396 => b:="5396";
                when 5397 => b:="5397";
                when 5398 => b:="5398";
                when 5399 => b:="5399";
                when 5400 => b:="5400";
                when 5401 => b:="5401";
                when 5402 => b:="5402";
                when 5403 => b:="5403";
                when 5404 => b:="5404";
                when 5405 => b:="5405";
                when 5406 => b:="5406";
                when 5407 => b:="5407";
                when 5408 => b:="5408";
                when 5409 => b:="5409";
                when 5410 => b:="5410";
                when 5411 => b:="5411";
                when 5412 => b:="5412";
                when 5413 => b:="5413";
                when 5414 => b:="5414";
                when 5415 => b:="5415";
                when 5416 => b:="5416";
                when 5417 => b:="5417";
                when 5418 => b:="5418";
                when 5419 => b:="5419";
                when 5420 => b:="5420";
                when 5421 => b:="5421";
                when 5422 => b:="5422";
                when 5423 => b:="5423";
                when 5424 => b:="5424";
                when 5425 => b:="5425";
                when 5426 => b:="5426";
                when 5427 => b:="5427";
                when 5428 => b:="5428";
                when 5429 => b:="5429";
                when 5430 => b:="5430";
                when 5431 => b:="5431";
                when 5432 => b:="5432";
                when 5433 => b:="5433";
                when 5434 => b:="5434";
                when 5435 => b:="5435";
                when 5436 => b:="5436";
                when 5437 => b:="5437";
                when 5438 => b:="5438";
                when 5439 => b:="5439";
                when 5440 => b:="5440";
                when 5441 => b:="5441";
                when 5442 => b:="5442";
                when 5443 => b:="5443";
                when 5444 => b:="5444";
                when 5445 => b:="5445";
                when 5446 => b:="5446";
                when 5447 => b:="5447";
                when 5448 => b:="5448";
                when 5449 => b:="5449";
                when 5450 => b:="5450";
                when 5451 => b:="5451";
                when 5452 => b:="5452";
                when 5453 => b:="5453";
                when 5454 => b:="5454";
                when 5455 => b:="5455";
                when 5456 => b:="5456";
                when 5457 => b:="5457";
                when 5458 => b:="5458";
                when 5459 => b:="5459";
                when 5460 => b:="5460";
                when 5461 => b:="5461";
                when 5462 => b:="5462";
                when 5463 => b:="5463";
                when 5464 => b:="5464";
                when 5465 => b:="5465";
                when 5466 => b:="5466";
                when 5467 => b:="5467";
                when 5468 => b:="5468";
                when 5469 => b:="5469";
                when 5470 => b:="5470";
                when 5471 => b:="5471";
                when 5472 => b:="5472";
                when 5473 => b:="5473";
                when 5474 => b:="5474";
                when 5475 => b:="5475";
                when 5476 => b:="5476";
                when 5477 => b:="5477";
                when 5478 => b:="5478";
                when 5479 => b:="5479";
                when 5480 => b:="5480";
                when 5481 => b:="5481";
                when 5482 => b:="5482";
                when 5483 => b:="5483";
                when 5484 => b:="5484";
                when 5485 => b:="5485";
                when 5486 => b:="5486";
                when 5487 => b:="5487";
                when 5488 => b:="5488";
                when 5489 => b:="5489";
                when 5490 => b:="5490";
                when 5491 => b:="5491";
                when 5492 => b:="5492";
                when 5493 => b:="5493";
                when 5494 => b:="5494";
                when 5495 => b:="5495";
                when 5496 => b:="5496";
                when 5497 => b:="5497";
                when 5498 => b:="5498";
                when 5499 => b:="5499";
                when 5500 => b:="5500";
                when 5501 => b:="5501";
                when 5502 => b:="5502";
                when 5503 => b:="5503";
                when 5504 => b:="5504";
                when 5505 => b:="5505";
                when 5506 => b:="5506";
                when 5507 => b:="5507";
                when 5508 => b:="5508";
                when 5509 => b:="5509";
                when 5510 => b:="5510";
                when 5511 => b:="5511";
                when 5512 => b:="5512";
                when 5513 => b:="5513";
                when 5514 => b:="5514";
                when 5515 => b:="5515";
                when 5516 => b:="5516";
                when 5517 => b:="5517";
                when 5518 => b:="5518";
                when 5519 => b:="5519";
                when 5520 => b:="5520";
                when 5521 => b:="5521";
                when 5522 => b:="5522";
                when 5523 => b:="5523";
                when 5524 => b:="5524";
                when 5525 => b:="5525";
                when 5526 => b:="5526";
                when 5527 => b:="5527";
                when 5528 => b:="5528";
                when 5529 => b:="5529";
                when 5530 => b:="5530";
                when 5531 => b:="5531";
                when 5532 => b:="5532";
                when 5533 => b:="5533";
                when 5534 => b:="5534";
                when 5535 => b:="5535";
                when 5536 => b:="5536";
                when 5537 => b:="5537";
                when 5538 => b:="5538";
                when 5539 => b:="5539";
                when 5540 => b:="5540";
                when 5541 => b:="5541";
                when 5542 => b:="5542";
                when 5543 => b:="5543";
                when 5544 => b:="5544";
                when 5545 => b:="5545";
                when 5546 => b:="5546";
                when 5547 => b:="5547";
                when 5548 => b:="5548";
                when 5549 => b:="5549";
                when 5550 => b:="5550";
                when 5551 => b:="5551";
                when 5552 => b:="5552";
                when 5553 => b:="5553";
                when 5554 => b:="5554";
                when 5555 => b:="5555";
                when 5556 => b:="5556";
                when 5557 => b:="5557";
                when 5558 => b:="5558";
                when 5559 => b:="5559";
                when 5560 => b:="5560";
                when 5561 => b:="5561";
                when 5562 => b:="5562";
                when 5563 => b:="5563";
                when 5564 => b:="5564";
                when 5565 => b:="5565";
                when 5566 => b:="5566";
                when 5567 => b:="5567";
                when 5568 => b:="5568";
                when 5569 => b:="5569";
                when 5570 => b:="5570";
                when 5571 => b:="5571";
                when 5572 => b:="5572";
                when 5573 => b:="5573";
                when 5574 => b:="5574";
                when 5575 => b:="5575";
                when 5576 => b:="5576";
                when 5577 => b:="5577";
                when 5578 => b:="5578";
                when 5579 => b:="5579";
                when 5580 => b:="5580";
                when 5581 => b:="5581";
                when 5582 => b:="5582";
                when 5583 => b:="5583";
                when 5584 => b:="5584";
                when 5585 => b:="5585";
                when 5586 => b:="5586";
                when 5587 => b:="5587";
                when 5588 => b:="5588";
                when 5589 => b:="5589";
                when 5590 => b:="5590";
                when 5591 => b:="5591";
                when 5592 => b:="5592";
                when 5593 => b:="5593";
                when 5594 => b:="5594";
                when 5595 => b:="5595";
                when 5596 => b:="5596";
                when 5597 => b:="5597";
                when 5598 => b:="5598";
                when 5599 => b:="5599";
                when 5600 => b:="5600";
                when 5601 => b:="5601";
                when 5602 => b:="5602";
                when 5603 => b:="5603";
                when 5604 => b:="5604";
                when 5605 => b:="5605";
                when 5606 => b:="5606";
                when 5607 => b:="5607";
                when 5608 => b:="5608";
                when 5609 => b:="5609";
                when 5610 => b:="5610";
                when 5611 => b:="5611";
                when 5612 => b:="5612";
                when 5613 => b:="5613";
                when 5614 => b:="5614";
                when 5615 => b:="5615";
                when 5616 => b:="5616";
                when 5617 => b:="5617";
                when 5618 => b:="5618";
                when 5619 => b:="5619";
                when 5620 => b:="5620";
                when 5621 => b:="5621";
                when 5622 => b:="5622";
                when 5623 => b:="5623";
                when 5624 => b:="5624";
                when 5625 => b:="5625";
                when 5626 => b:="5626";
                when 5627 => b:="5627";
                when 5628 => b:="5628";
                when 5629 => b:="5629";
                when 5630 => b:="5630";
                when 5631 => b:="5631";
                when 5632 => b:="5632";
                when 5633 => b:="5633";
                when 5634 => b:="5634";
                when 5635 => b:="5635";
                when 5636 => b:="5636";
                when 5637 => b:="5637";
                when 5638 => b:="5638";
                when 5639 => b:="5639";
                when 5640 => b:="5640";
                when 5641 => b:="5641";
                when 5642 => b:="5642";
                when 5643 => b:="5643";
                when 5644 => b:="5644";
                when 5645 => b:="5645";
                when 5646 => b:="5646";
                when 5647 => b:="5647";
                when 5648 => b:="5648";
                when 5649 => b:="5649";
                when 5650 => b:="5650";
                when 5651 => b:="5651";
                when 5652 => b:="5652";
                when 5653 => b:="5653";
                when 5654 => b:="5654";
                when 5655 => b:="5655";
                when 5656 => b:="5656";
                when 5657 => b:="5657";
                when 5658 => b:="5658";
                when 5659 => b:="5659";
                when 5660 => b:="5660";
                when 5661 => b:="5661";
                when 5662 => b:="5662";
                when 5663 => b:="5663";
                when 5664 => b:="5664";
                when 5665 => b:="5665";
                when 5666 => b:="5666";
                when 5667 => b:="5667";
                when 5668 => b:="5668";
                when 5669 => b:="5669";
                when 5670 => b:="5670";
                when 5671 => b:="5671";
                when 5672 => b:="5672";
                when 5673 => b:="5673";
                when 5674 => b:="5674";
                when 5675 => b:="5675";
                when 5676 => b:="5676";
                when 5677 => b:="5677";
                when 5678 => b:="5678";
                when 5679 => b:="5679";
                when 5680 => b:="5680";
                when 5681 => b:="5681";
                when 5682 => b:="5682";
                when 5683 => b:="5683";
                when 5684 => b:="5684";
                when 5685 => b:="5685";
                when 5686 => b:="5686";
                when 5687 => b:="5687";
                when 5688 => b:="5688";
                when 5689 => b:="5689";
                when 5690 => b:="5690";
                when 5691 => b:="5691";
                when 5692 => b:="5692";
                when 5693 => b:="5693";
                when 5694 => b:="5694";
                when 5695 => b:="5695";
                when 5696 => b:="5696";
                when 5697 => b:="5697";
                when 5698 => b:="5698";
                when 5699 => b:="5699";
                when 5700 => b:="5700";
                when 5701 => b:="5701";
                when 5702 => b:="5702";
                when 5703 => b:="5703";
                when 5704 => b:="5704";
                when 5705 => b:="5705";
                when 5706 => b:="5706";
                when 5707 => b:="5707";
                when 5708 => b:="5708";
                when 5709 => b:="5709";
                when 5710 => b:="5710";
                when 5711 => b:="5711";
                when 5712 => b:="5712";
                when 5713 => b:="5713";
                when 5714 => b:="5714";
                when 5715 => b:="5715";
                when 5716 => b:="5716";
                when 5717 => b:="5717";
                when 5718 => b:="5718";
                when 5719 => b:="5719";
                when 5720 => b:="5720";
                when 5721 => b:="5721";
                when 5722 => b:="5722";
                when 5723 => b:="5723";
                when 5724 => b:="5724";
                when 5725 => b:="5725";
                when 5726 => b:="5726";
                when 5727 => b:="5727";
                when 5728 => b:="5728";
                when 5729 => b:="5729";
                when 5730 => b:="5730";
                when 5731 => b:="5731";
                when 5732 => b:="5732";
                when 5733 => b:="5733";
                when 5734 => b:="5734";
                when 5735 => b:="5735";
                when 5736 => b:="5736";
                when 5737 => b:="5737";
                when 5738 => b:="5738";
                when 5739 => b:="5739";
                when 5740 => b:="5740";
                when 5741 => b:="5741";
                when 5742 => b:="5742";
                when 5743 => b:="5743";
                when 5744 => b:="5744";
                when 5745 => b:="5745";
                when 5746 => b:="5746";
                when 5747 => b:="5747";
                when 5748 => b:="5748";
                when 5749 => b:="5749";
                when 5750 => b:="5750";
                when 5751 => b:="5751";
                when 5752 => b:="5752";
                when 5753 => b:="5753";
                when 5754 => b:="5754";
                when 5755 => b:="5755";
                when 5756 => b:="5756";
                when 5757 => b:="5757";
                when 5758 => b:="5758";
                when 5759 => b:="5759";
                when 5760 => b:="5760";
                when 5761 => b:="5761";
                when 5762 => b:="5762";
                when 5763 => b:="5763";
                when 5764 => b:="5764";
                when 5765 => b:="5765";
                when 5766 => b:="5766";
                when 5767 => b:="5767";
                when 5768 => b:="5768";
                when 5769 => b:="5769";
                when 5770 => b:="5770";
                when 5771 => b:="5771";
                when 5772 => b:="5772";
                when 5773 => b:="5773";
                when 5774 => b:="5774";
                when 5775 => b:="5775";
                when 5776 => b:="5776";
                when 5777 => b:="5777";
                when 5778 => b:="5778";
                when 5779 => b:="5779";
                when 5780 => b:="5780";
                when 5781 => b:="5781";
                when 5782 => b:="5782";
                when 5783 => b:="5783";
                when 5784 => b:="5784";
                when 5785 => b:="5785";
                when 5786 => b:="5786";
                when 5787 => b:="5787";
                when 5788 => b:="5788";
                when 5789 => b:="5789";
                when 5790 => b:="5790";
                when 5791 => b:="5791";
                when 5792 => b:="5792";
                when 5793 => b:="5793";
                when 5794 => b:="5794";
                when 5795 => b:="5795";
                when 5796 => b:="5796";
                when 5797 => b:="5797";
                when 5798 => b:="5798";
                when 5799 => b:="5799";
                when 5800 => b:="5800";
                when 5801 => b:="5801";
                when 5802 => b:="5802";
                when 5803 => b:="5803";
                when 5804 => b:="5804";
                when 5805 => b:="5805";
                when 5806 => b:="5806";
                when 5807 => b:="5807";
                when 5808 => b:="5808";
                when 5809 => b:="5809";
                when 5810 => b:="5810";
                when 5811 => b:="5811";
                when 5812 => b:="5812";
                when 5813 => b:="5813";
                when 5814 => b:="5814";
                when 5815 => b:="5815";
                when 5816 => b:="5816";
                when 5817 => b:="5817";
                when 5818 => b:="5818";
                when 5819 => b:="5819";
                when 5820 => b:="5820";
                when 5821 => b:="5821";
                when 5822 => b:="5822";
                when 5823 => b:="5823";
                when 5824 => b:="5824";
                when 5825 => b:="5825";
                when 5826 => b:="5826";
                when 5827 => b:="5827";
                when 5828 => b:="5828";
                when 5829 => b:="5829";
                when 5830 => b:="5830";
                when 5831 => b:="5831";
                when 5832 => b:="5832";
                when 5833 => b:="5833";
                when 5834 => b:="5834";
                when 5835 => b:="5835";
                when 5836 => b:="5836";
                when 5837 => b:="5837";
                when 5838 => b:="5838";
                when 5839 => b:="5839";
                when 5840 => b:="5840";
                when 5841 => b:="5841";
                when 5842 => b:="5842";
                when 5843 => b:="5843";
                when 5844 => b:="5844";
                when 5845 => b:="5845";
                when 5846 => b:="5846";
                when 5847 => b:="5847";
                when 5848 => b:="5848";
                when 5849 => b:="5849";
                when 5850 => b:="5850";
                when 5851 => b:="5851";
                when 5852 => b:="5852";
                when 5853 => b:="5853";
                when 5854 => b:="5854";
                when 5855 => b:="5855";
                when 5856 => b:="5856";
                when 5857 => b:="5857";
                when 5858 => b:="5858";
                when 5859 => b:="5859";
                when 5860 => b:="5860";
                when 5861 => b:="5861";
                when 5862 => b:="5862";
                when 5863 => b:="5863";
                when 5864 => b:="5864";
                when 5865 => b:="5865";
                when 5866 => b:="5866";
                when 5867 => b:="5867";
                when 5868 => b:="5868";
                when 5869 => b:="5869";
                when 5870 => b:="5870";
                when 5871 => b:="5871";
                when 5872 => b:="5872";
                when 5873 => b:="5873";
                when 5874 => b:="5874";
                when 5875 => b:="5875";
                when 5876 => b:="5876";
                when 5877 => b:="5877";
                when 5878 => b:="5878";
                when 5879 => b:="5879";
                when 5880 => b:="5880";
                when 5881 => b:="5881";
                when 5882 => b:="5882";
                when 5883 => b:="5883";
                when 5884 => b:="5884";
                when 5885 => b:="5885";
                when 5886 => b:="5886";
                when 5887 => b:="5887";
                when 5888 => b:="5888";
                when 5889 => b:="5889";
                when 5890 => b:="5890";
                when 5891 => b:="5891";
                when 5892 => b:="5892";
                when 5893 => b:="5893";
                when 5894 => b:="5894";
                when 5895 => b:="5895";
                when 5896 => b:="5896";
                when 5897 => b:="5897";
                when 5898 => b:="5898";
                when 5899 => b:="5899";
                when 5900 => b:="5900";
                when 5901 => b:="5901";
                when 5902 => b:="5902";
                when 5903 => b:="5903";
                when 5904 => b:="5904";
                when 5905 => b:="5905";
                when 5906 => b:="5906";
                when 5907 => b:="5907";
                when 5908 => b:="5908";
                when 5909 => b:="5909";
                when 5910 => b:="5910";
                when 5911 => b:="5911";
                when 5912 => b:="5912";
                when 5913 => b:="5913";
                when 5914 => b:="5914";
                when 5915 => b:="5915";
                when 5916 => b:="5916";
                when 5917 => b:="5917";
                when 5918 => b:="5918";
                when 5919 => b:="5919";
                when 5920 => b:="5920";
                when 5921 => b:="5921";
                when 5922 => b:="5922";
                when 5923 => b:="5923";
                when 5924 => b:="5924";
                when 5925 => b:="5925";
                when 5926 => b:="5926";
                when 5927 => b:="5927";
                when 5928 => b:="5928";
                when 5929 => b:="5929";
                when 5930 => b:="5930";
                when 5931 => b:="5931";
                when 5932 => b:="5932";
                when 5933 => b:="5933";
                when 5934 => b:="5934";
                when 5935 => b:="5935";
                when 5936 => b:="5936";
                when 5937 => b:="5937";
                when 5938 => b:="5938";
                when 5939 => b:="5939";
                when 5940 => b:="5940";
                when 5941 => b:="5941";
                when 5942 => b:="5942";
                when 5943 => b:="5943";
                when 5944 => b:="5944";
                when 5945 => b:="5945";
                when 5946 => b:="5946";
                when 5947 => b:="5947";
                when 5948 => b:="5948";
                when 5949 => b:="5949";
                when 5950 => b:="5950";
                when 5951 => b:="5951";
                when 5952 => b:="5952";
                when 5953 => b:="5953";
                when 5954 => b:="5954";
                when 5955 => b:="5955";
                when 5956 => b:="5956";
                when 5957 => b:="5957";
                when 5958 => b:="5958";
                when 5959 => b:="5959";
                when 5960 => b:="5960";
                when 5961 => b:="5961";
                when 5962 => b:="5962";
                when 5963 => b:="5963";
                when 5964 => b:="5964";
                when 5965 => b:="5965";
                when 5966 => b:="5966";
                when 5967 => b:="5967";
                when 5968 => b:="5968";
                when 5969 => b:="5969";
                when 5970 => b:="5970";
                when 5971 => b:="5971";
                when 5972 => b:="5972";
                when 5973 => b:="5973";
                when 5974 => b:="5974";
                when 5975 => b:="5975";
                when 5976 => b:="5976";
                when 5977 => b:="5977";
                when 5978 => b:="5978";
                when 5979 => b:="5979";
                when 5980 => b:="5980";
                when 5981 => b:="5981";
                when 5982 => b:="5982";
                when 5983 => b:="5983";
                when 5984 => b:="5984";
                when 5985 => b:="5985";
                when 5986 => b:="5986";
                when 5987 => b:="5987";
                when 5988 => b:="5988";
                when 5989 => b:="5989";
                when 5990 => b:="5990";
                when 5991 => b:="5991";
                when 5992 => b:="5992";
                when 5993 => b:="5993";
                when 5994 => b:="5994";
                when 5995 => b:="5995";
                when 5996 => b:="5996";
                when 5997 => b:="5997";
                when 5998 => b:="5998";
                when 6000 => b:="6000";
                when 6001 => b:="6001";
                when 6002 => b:="6002";
                when 6003 => b:="6003";
                when 6004 => b:="6004";
                when 6005 => b:="6005";
                when 6006 => b:="6006";
                when 6007 => b:="6007";
                when 6008 => b:="6008";
                when 6009 => b:="6009";
                when 6010 => b:="6010";
                when 6011 => b:="6011";
                when 6012 => b:="6012";
                when 6013 => b:="6013";
                when 6014 => b:="6014";
                when 6015 => b:="6015";
                when 6016 => b:="6016";
                when 6017 => b:="6017";
                when 6018 => b:="6018";
                when 6019 => b:="6019";
                when 6020 => b:="6020";
                when 6021 => b:="6021";
                when 6022 => b:="6022";
                when 6023 => b:="6023";
                when 6024 => b:="6024";
                when 6025 => b:="6025";
                when 6026 => b:="6026";
                when 6027 => b:="6027";
                when 6028 => b:="6028";
                when 6029 => b:="6029";
                when 6030 => b:="6030";
                when 6031 => b:="6031";
                when 6032 => b:="6032";
                when 6033 => b:="6033";
                when 6034 => b:="6034";
                when 6035 => b:="6035";
                when 6036 => b:="6036";
                when 6037 => b:="6037";
                when 6038 => b:="6038";
                when 6039 => b:="6039";
                when 6040 => b:="6040";
                when 6041 => b:="6041";
                when 6042 => b:="6042";
                when 6043 => b:="6043";
                when 6044 => b:="6044";
                when 6045 => b:="6045";
                when 6046 => b:="6046";
                when 6047 => b:="6047";
                when 6048 => b:="6048";
                when 6049 => b:="6049";
                when 6050 => b:="6050";
                when 6051 => b:="6051";
                when 6052 => b:="6052";
                when 6053 => b:="6053";
                when 6054 => b:="6054";
                when 6055 => b:="6055";
                when 6056 => b:="6056";
                when 6057 => b:="6057";
                when 6058 => b:="6058";
                when 6059 => b:="6059";
                when 6060 => b:="6060";
                when 6061 => b:="6061";
                when 6062 => b:="6062";
                when 6063 => b:="6063";
                when 6064 => b:="6064";
                when 6065 => b:="6065";
                when 6066 => b:="6066";
                when 6067 => b:="6067";
                when 6068 => b:="6068";
                when 6069 => b:="6069";
                when 6070 => b:="6070";
                when 6071 => b:="6071";
                when 6072 => b:="6072";
                when 6073 => b:="6073";
                when 6074 => b:="6074";
                when 6075 => b:="6075";
                when 6076 => b:="6076";
                when 6077 => b:="6077";
                when 6078 => b:="6078";
                when 6079 => b:="6079";
                when 6080 => b:="6080";
                when 6081 => b:="6081";
                when 6082 => b:="6082";
                when 6083 => b:="6083";
                when 6084 => b:="6084";
                when 6085 => b:="6085";
                when 6086 => b:="6086";
                when 6087 => b:="6087";
                when 6088 => b:="6088";
                when 6089 => b:="6089";
                when 6090 => b:="6090";
                when 6091 => b:="6091";
                when 6092 => b:="6092";
                when 6093 => b:="6093";
                when 6094 => b:="6094";
                when 6095 => b:="6095";
                when 6096 => b:="6096";
                when 6097 => b:="6097";
                when 6098 => b:="6098";
                when 6099 => b:="6099";
                when 6100 => b:="6100";
                when 6101 => b:="6101";
                when 6102 => b:="6102";
                when 6103 => b:="6103";
                when 6104 => b:="6104";
                when 6105 => b:="6105";
                when 6106 => b:="6106";
                when 6107 => b:="6107";
                when 6108 => b:="6108";
                when 6109 => b:="6109";
                when 6110 => b:="6110";
                when 6111 => b:="6111";
                when 6112 => b:="6112";
                when 6113 => b:="6113";
                when 6114 => b:="6114";
                when 6115 => b:="6115";
                when 6116 => b:="6116";
                when 6117 => b:="6117";
                when 6118 => b:="6118";
                when 6119 => b:="6119";
                when 6120 => b:="6120";
                when 6121 => b:="6121";
                when 6122 => b:="6122";
                when 6123 => b:="6123";
                when 6124 => b:="6124";
                when 6125 => b:="6125";
                when 6126 => b:="6126";
                when 6127 => b:="6127";
                when 6128 => b:="6128";
                when 6129 => b:="6129";
                when 6130 => b:="6130";
                when 6131 => b:="6131";
                when 6132 => b:="6132";
                when 6133 => b:="6133";
                when 6134 => b:="6134";
                when 6135 => b:="6135";
                when 6136 => b:="6136";
                when 6137 => b:="6137";
                when 6138 => b:="6138";
                when 6139 => b:="6139";
                when 6140 => b:="6140";
                when 6141 => b:="6141";
                when 6142 => b:="6142";
                when 6143 => b:="6143";
                when 6144 => b:="6144";
                when 6145 => b:="6145";
                when 6146 => b:="6146";
                when 6147 => b:="6147";
                when 6148 => b:="6148";
                when 6149 => b:="6149";
                when 6150 => b:="6150";
                when 6151 => b:="6151";
                when 6152 => b:="6152";
                when 6153 => b:="6153";
                when 6154 => b:="6154";
                when 6155 => b:="6155";
                when 6156 => b:="6156";
                when 6157 => b:="6157";
                when 6158 => b:="6158";
                when 6159 => b:="6159";
                when 6160 => b:="6160";
                when 6161 => b:="6161";
                when 6162 => b:="6162";
                when 6163 => b:="6163";
                when 6164 => b:="6164";
                when 6165 => b:="6165";
                when 6166 => b:="6166";
                when 6167 => b:="6167";
                when 6168 => b:="6168";
                when 6169 => b:="6169";
                when 6170 => b:="6170";
                when 6171 => b:="6171";
                when 6172 => b:="6172";
                when 6173 => b:="6173";
                when 6174 => b:="6174";
                when 6175 => b:="6175";
                when 6176 => b:="6176";
                when 6177 => b:="6177";
                when 6178 => b:="6178";
                when 6179 => b:="6179";
                when 6180 => b:="6180";
                when 6181 => b:="6181";
                when 6182 => b:="6182";
                when 6183 => b:="6183";
                when 6184 => b:="6184";
                when 6185 => b:="6185";
                when 6186 => b:="6186";
                when 6187 => b:="6187";
                when 6188 => b:="6188";
                when 6189 => b:="6189";
                when 6190 => b:="6190";
                when 6191 => b:="6191";
                when 6192 => b:="6192";
                when 6193 => b:="6193";
                when 6194 => b:="6194";
                when 6195 => b:="6195";
                when 6196 => b:="6196";
                when 6197 => b:="6197";
                when 6198 => b:="6198";
                when 6199 => b:="6199";
                when 6200 => b:="6200";
                when 6201 => b:="6201";
                when 6202 => b:="6202";
                when 6203 => b:="6203";
                when 6204 => b:="6204";
                when 6205 => b:="6205";
                when 6206 => b:="6206";
                when 6207 => b:="6207";
                when 6208 => b:="6208";
                when 6209 => b:="6209";
                when 6210 => b:="6210";
                when 6211 => b:="6211";
                when 6212 => b:="6212";
                when 6213 => b:="6213";
                when 6214 => b:="6214";
                when 6215 => b:="6215";
                when 6216 => b:="6216";
                when 6217 => b:="6217";
                when 6218 => b:="6218";
                when 6219 => b:="6219";
                when 6220 => b:="6220";
                when 6221 => b:="6221";
                when 6222 => b:="6222";
                when 6223 => b:="6223";
                when 6224 => b:="6224";
                when 6225 => b:="6225";
                when 6226 => b:="6226";
                when 6227 => b:="6227";
                when 6228 => b:="6228";
                when 6229 => b:="6229";
                when 6230 => b:="6230";
                when 6231 => b:="6231";
                when 6232 => b:="6232";
                when 6233 => b:="6233";
                when 6234 => b:="6234";
                when 6235 => b:="6235";
                when 6236 => b:="6236";
                when 6237 => b:="6237";
                when 6238 => b:="6238";
                when 6239 => b:="6239";
                when 6240 => b:="6240";
                when 6241 => b:="6241";
                when 6242 => b:="6242";
                when 6243 => b:="6243";
                when 6244 => b:="6244";
                when 6245 => b:="6245";
                when 6246 => b:="6246";
                when 6247 => b:="6247";
                when 6248 => b:="6248";
                when 6249 => b:="6249";
                when 6250 => b:="6250";
                when 6251 => b:="6251";
                when 6252 => b:="6252";
                when 6253 => b:="6253";
                when 6254 => b:="6254";
                when 6255 => b:="6255";
                when 6256 => b:="6256";
                when 6257 => b:="6257";
                when 6258 => b:="6258";
                when 6259 => b:="6259";
                when 6260 => b:="6260";
                when 6261 => b:="6261";
                when 6262 => b:="6262";
                when 6263 => b:="6263";
                when 6264 => b:="6264";
                when 6265 => b:="6265";
                when 6266 => b:="6266";
                when 6267 => b:="6267";
                when 6268 => b:="6268";
                when 6269 => b:="6269";
                when 6270 => b:="6270";
                when 6271 => b:="6271";
                when 6272 => b:="6272";
                when 6273 => b:="6273";
                when 6274 => b:="6274";
                when 6275 => b:="6275";
                when 6276 => b:="6276";
                when 6277 => b:="6277";
                when 6278 => b:="6278";
                when 6279 => b:="6279";
                when 6280 => b:="6280";
                when 6281 => b:="6281";
                when 6282 => b:="6282";
                when 6283 => b:="6283";
                when 6284 => b:="6284";
                when 6285 => b:="6285";
                when 6286 => b:="6286";
                when 6287 => b:="6287";
                when 6288 => b:="6288";
                when 6289 => b:="6289";
                when 6290 => b:="6290";
                when 6291 => b:="6291";
                when 6292 => b:="6292";
                when 6293 => b:="6293";
                when 6294 => b:="6294";
                when 6295 => b:="6295";
                when 6296 => b:="6296";
                when 6297 => b:="6297";
                when 6298 => b:="6298";
                when 6299 => b:="6299";
                when 6300 => b:="6300";
                when 6301 => b:="6301";
                when 6302 => b:="6302";
                when 6303 => b:="6303";
                when 6304 => b:="6304";
                when 6305 => b:="6305";
                when 6306 => b:="6306";
                when 6307 => b:="6307";
                when 6308 => b:="6308";
                when 6309 => b:="6309";
                when 6310 => b:="6310";
                when 6311 => b:="6311";
                when 6312 => b:="6312";
                when 6313 => b:="6313";
                when 6314 => b:="6314";
                when 6315 => b:="6315";
                when 6316 => b:="6316";
                when 6317 => b:="6317";
                when 6318 => b:="6318";
                when 6319 => b:="6319";
                when 6320 => b:="6320";
                when 6321 => b:="6321";
                when 6322 => b:="6322";
                when 6323 => b:="6323";
                when 6324 => b:="6324";
                when 6325 => b:="6325";
                when 6326 => b:="6326";
                when 6327 => b:="6327";
                when 6328 => b:="6328";
                when 6329 => b:="6329";
                when 6330 => b:="6330";
                when 6331 => b:="6331";
                when 6332 => b:="6332";
                when 6333 => b:="6333";
                when 6334 => b:="6334";
                when 6335 => b:="6335";
                when 6336 => b:="6336";
                when 6337 => b:="6337";
                when 6338 => b:="6338";
                when 6339 => b:="6339";
                when 6340 => b:="6340";
                when 6341 => b:="6341";
                when 6342 => b:="6342";
                when 6343 => b:="6343";
                when 6344 => b:="6344";
                when 6345 => b:="6345";
                when 6346 => b:="6346";
                when 6347 => b:="6347";
                when 6348 => b:="6348";
                when 6349 => b:="6349";
                when 6350 => b:="6350";
                when 6351 => b:="6351";
                when 6352 => b:="6352";
                when 6353 => b:="6353";
                when 6354 => b:="6354";
                when 6355 => b:="6355";
                when 6356 => b:="6356";
                when 6357 => b:="6357";
                when 6358 => b:="6358";
                when 6359 => b:="6359";
                when 6360 => b:="6360";
                when 6361 => b:="6361";
                when 6362 => b:="6362";
                when 6363 => b:="6363";
                when 6364 => b:="6364";
                when 6365 => b:="6365";
                when 6366 => b:="6366";
                when 6367 => b:="6367";
                when 6368 => b:="6368";
                when 6369 => b:="6369";
                when 6370 => b:="6370";
                when 6371 => b:="6371";
                when 6372 => b:="6372";
                when 6373 => b:="6373";
                when 6374 => b:="6374";
                when 6375 => b:="6375";
                when 6376 => b:="6376";
                when 6377 => b:="6377";
                when 6378 => b:="6378";
                when 6379 => b:="6379";
                when 6380 => b:="6380";
                when 6381 => b:="6381";
                when 6382 => b:="6382";
                when 6383 => b:="6383";
                when 6384 => b:="6384";
                when 6385 => b:="6385";
                when 6386 => b:="6386";
                when 6387 => b:="6387";
                when 6388 => b:="6388";
                when 6389 => b:="6389";
                when 6390 => b:="6390";
                when 6391 => b:="6391";
                when 6392 => b:="6392";
                when 6393 => b:="6393";
                when 6394 => b:="6394";
                when 6395 => b:="6395";
                when 6396 => b:="6396";
                when 6397 => b:="6397";
                when 6398 => b:="6398";
                when 6399 => b:="6399";
                when 6400 => b:="6400";
                when 6401 => b:="6401";
                when 6402 => b:="6402";
                when 6403 => b:="6403";
                when 6404 => b:="6404";
                when 6405 => b:="6405";
                when 6406 => b:="6406";
                when 6407 => b:="6407";
                when 6408 => b:="6408";
                when 6409 => b:="6409";
                when 6410 => b:="6410";
                when 6411 => b:="6411";
                when 6412 => b:="6412";
                when 6413 => b:="6413";
                when 6414 => b:="6414";
                when 6415 => b:="6415";
                when 6416 => b:="6416";
                when 6417 => b:="6417";
                when 6418 => b:="6418";
                when 6419 => b:="6419";
                when 6420 => b:="6420";
                when 6421 => b:="6421";
                when 6422 => b:="6422";
                when 6423 => b:="6423";
                when 6424 => b:="6424";
                when 6425 => b:="6425";
                when 6426 => b:="6426";
                when 6427 => b:="6427";
                when 6428 => b:="6428";
                when 6429 => b:="6429";
                when 6430 => b:="6430";
                when 6431 => b:="6431";
                when 6432 => b:="6432";
                when 6433 => b:="6433";
                when 6434 => b:="6434";
                when 6435 => b:="6435";
                when 6436 => b:="6436";
                when 6437 => b:="6437";
                when 6438 => b:="6438";
                when 6439 => b:="6439";
                when 6440 => b:="6440";
                when 6441 => b:="6441";
                when 6442 => b:="6442";
                when 6443 => b:="6443";
                when 6444 => b:="6444";
                when 6445 => b:="6445";
                when 6446 => b:="6446";
                when 6447 => b:="6447";
                when 6448 => b:="6448";
                when 6449 => b:="6449";
                when 6450 => b:="6450";
                when 6451 => b:="6451";
                when 6452 => b:="6452";
                when 6453 => b:="6453";
                when 6454 => b:="6454";
                when 6455 => b:="6455";
                when 6456 => b:="6456";
                when 6457 => b:="6457";
                when 6458 => b:="6458";
                when 6459 => b:="6459";
                when 6460 => b:="6460";
                when 6461 => b:="6461";
                when 6462 => b:="6462";
                when 6463 => b:="6463";
                when 6464 => b:="6464";
                when 6465 => b:="6465";
                when 6466 => b:="6466";
                when 6467 => b:="6467";
                when 6468 => b:="6468";
                when 6469 => b:="6469";
                when 6470 => b:="6470";
                when 6471 => b:="6471";
                when 6472 => b:="6472";
                when 6473 => b:="6473";
                when 6474 => b:="6474";
                when 6475 => b:="6475";
                when 6476 => b:="6476";
                when 6477 => b:="6477";
                when 6478 => b:="6478";
                when 6479 => b:="6479";
                when 6480 => b:="6480";
                when 6481 => b:="6481";
                when 6482 => b:="6482";
                when 6483 => b:="6483";
                when 6484 => b:="6484";
                when 6485 => b:="6485";
                when 6486 => b:="6486";
                when 6487 => b:="6487";
                when 6488 => b:="6488";
                when 6489 => b:="6489";
                when 6490 => b:="6490";
                when 6491 => b:="6491";
                when 6492 => b:="6492";
                when 6493 => b:="6493";
                when 6494 => b:="6494";
                when 6495 => b:="6495";
                when 6496 => b:="6496";
                when 6497 => b:="6497";
                when 6498 => b:="6498";
                when 6499 => b:="6499";
                when 6500 => b:="6500";
                when 6501 => b:="6501";
                when 6502 => b:="6502";
                when 6503 => b:="6503";
                when 6504 => b:="6504";
                when 6505 => b:="6505";
                when 6506 => b:="6506";
                when 6507 => b:="6507";
                when 6508 => b:="6508";
                when 6509 => b:="6509";
                when 6510 => b:="6510";
                when 6511 => b:="6511";
                when 6512 => b:="6512";
                when 6513 => b:="6513";
                when 6514 => b:="6514";
                when 6515 => b:="6515";
                when 6516 => b:="6516";
                when 6517 => b:="6517";
                when 6518 => b:="6518";
                when 6519 => b:="6519";
                when 6520 => b:="6520";
                when 6521 => b:="6521";
                when 6522 => b:="6522";
                when 6523 => b:="6523";
                when 6524 => b:="6524";
                when 6525 => b:="6525";
                when 6526 => b:="6526";
                when 6527 => b:="6527";
                when 6528 => b:="6528";
                when 6529 => b:="6529";
                when 6530 => b:="6530";
                when 6531 => b:="6531";
                when 6532 => b:="6532";
                when 6533 => b:="6533";
                when 6534 => b:="6534";
                when 6535 => b:="6535";
                when 6536 => b:="6536";
                when 6537 => b:="6537";
                when 6538 => b:="6538";
                when 6539 => b:="6539";
                when 6540 => b:="6540";
                when 6541 => b:="6541";
                when 6542 => b:="6542";
                when 6543 => b:="6543";
                when 6544 => b:="6544";
                when 6545 => b:="6545";
                when 6546 => b:="6546";
                when 6547 => b:="6547";
                when 6548 => b:="6548";
                when 6549 => b:="6549";
                when 6550 => b:="6550";
                when 6551 => b:="6551";
                when 6552 => b:="6552";
                when 6553 => b:="6553";
                when 6554 => b:="6554";
                when 6555 => b:="6555";
                when 6556 => b:="6556";
                when 6557 => b:="6557";
                when 6558 => b:="6558";
                when 6559 => b:="6559";
                when 6560 => b:="6560";
                when 6561 => b:="6561";
                when 6562 => b:="6562";
                when 6563 => b:="6563";
                when 6564 => b:="6564";
                when 6565 => b:="6565";
                when 6566 => b:="6566";
                when 6567 => b:="6567";
                when 6568 => b:="6568";
                when 6569 => b:="6569";
                when 6570 => b:="6570";
                when 6571 => b:="6571";
                when 6572 => b:="6572";
                when 6573 => b:="6573";
                when 6574 => b:="6574";
                when 6575 => b:="6575";
                when 6576 => b:="6576";
                when 6577 => b:="6577";
                when 6578 => b:="6578";
                when 6579 => b:="6579";
                when 6580 => b:="6580";
                when 6581 => b:="6581";
                when 6582 => b:="6582";
                when 6583 => b:="6583";
                when 6584 => b:="6584";
                when 6585 => b:="6585";
                when 6586 => b:="6586";
                when 6587 => b:="6587";
                when 6588 => b:="6588";
                when 6589 => b:="6589";
                when 6590 => b:="6590";
                when 6591 => b:="6591";
                when 6592 => b:="6592";
                when 6593 => b:="6593";
                when 6594 => b:="6594";
                when 6595 => b:="6595";
                when 6596 => b:="6596";
                when 6597 => b:="6597";
                when 6598 => b:="6598";
                when 6599 => b:="6599";
                when 6600 => b:="6600";
                when 6601 => b:="6601";
                when 6602 => b:="6602";
                when 6603 => b:="6603";
                when 6604 => b:="6604";
                when 6605 => b:="6605";
                when 6606 => b:="6606";
                when 6607 => b:="6607";
                when 6608 => b:="6608";
                when 6609 => b:="6609";
                when 6610 => b:="6610";
                when 6611 => b:="6611";
                when 6612 => b:="6612";
                when 6613 => b:="6613";
                when 6614 => b:="6614";
                when 6615 => b:="6615";
                when 6616 => b:="6616";
                when 6617 => b:="6617";
                when 6618 => b:="6618";
                when 6619 => b:="6619";
                when 6620 => b:="6620";
                when 6621 => b:="6621";
                when 6622 => b:="6622";
                when 6623 => b:="6623";
                when 6624 => b:="6624";
                when 6625 => b:="6625";
                when 6626 => b:="6626";
                when 6627 => b:="6627";
                when 6628 => b:="6628";
                when 6629 => b:="6629";
                when 6630 => b:="6630";
                when 6631 => b:="6631";
                when 6632 => b:="6632";
                when 6633 => b:="6633";
                when 6634 => b:="6634";
                when 6635 => b:="6635";
                when 6636 => b:="6636";
                when 6637 => b:="6637";
                when 6638 => b:="6638";
                when 6639 => b:="6639";
                when 6640 => b:="6640";
                when 6641 => b:="6641";
                when 6642 => b:="6642";
                when 6643 => b:="6643";
                when 6644 => b:="6644";
                when 6645 => b:="6645";
                when 6646 => b:="6646";
                when 6647 => b:="6647";
                when 6648 => b:="6648";
                when 6649 => b:="6649";
                when 6650 => b:="6650";
                when 6651 => b:="6651";
                when 6652 => b:="6652";
                when 6653 => b:="6653";
                when 6654 => b:="6654";
                when 6655 => b:="6655";
                when 6656 => b:="6656";
                when 6657 => b:="6657";
                when 6658 => b:="6658";
                when 6659 => b:="6659";
                when 6660 => b:="6660";
                when 6661 => b:="6661";
                when 6662 => b:="6662";
                when 6663 => b:="6663";
                when 6664 => b:="6664";
                when 6665 => b:="6665";
                when 6666 => b:="6666";
                when 6667 => b:="6667";
                when 6668 => b:="6668";
                when 6669 => b:="6669";
                when 6670 => b:="6670";
                when 6671 => b:="6671";
                when 6672 => b:="6672";
                when 6673 => b:="6673";
                when 6674 => b:="6674";
                when 6675 => b:="6675";
                when 6676 => b:="6676";
                when 6677 => b:="6677";
                when 6678 => b:="6678";
                when 6679 => b:="6679";
                when 6680 => b:="6680";
                when 6681 => b:="6681";
                when 6682 => b:="6682";
                when 6683 => b:="6683";
                when 6684 => b:="6684";
                when 6685 => b:="6685";
                when 6686 => b:="6686";
                when 6687 => b:="6687";
                when 6688 => b:="6688";
                when 6689 => b:="6689";
                when 6690 => b:="6690";
                when 6691 => b:="6691";
                when 6692 => b:="6692";
                when 6693 => b:="6693";
                when 6694 => b:="6694";
                when 6695 => b:="6695";
                when 6696 => b:="6696";
                when 6697 => b:="6697";
                when 6698 => b:="6698";
                when 6699 => b:="6699";
                when 6700 => b:="6700";
                when 6701 => b:="6701";
                when 6702 => b:="6702";
                when 6703 => b:="6703";
                when 6704 => b:="6704";
                when 6705 => b:="6705";
                when 6706 => b:="6706";
                when 6707 => b:="6707";
                when 6708 => b:="6708";
                when 6709 => b:="6709";
                when 6710 => b:="6710";
                when 6711 => b:="6711";
                when 6712 => b:="6712";
                when 6713 => b:="6713";
                when 6714 => b:="6714";
                when 6715 => b:="6715";
                when 6716 => b:="6716";
                when 6717 => b:="6717";
                when 6718 => b:="6718";
                when 6719 => b:="6719";
                when 6720 => b:="6720";
                when 6721 => b:="6721";
                when 6722 => b:="6722";
                when 6723 => b:="6723";
                when 6724 => b:="6724";
                when 6725 => b:="6725";
                when 6726 => b:="6726";
                when 6727 => b:="6727";
                when 6728 => b:="6728";
                when 6729 => b:="6729";
                when 6730 => b:="6730";
                when 6731 => b:="6731";
                when 6732 => b:="6732";
                when 6733 => b:="6733";
                when 6734 => b:="6734";
                when 6735 => b:="6735";
                when 6736 => b:="6736";
                when 6737 => b:="6737";
                when 6738 => b:="6738";
                when 6739 => b:="6739";
                when 6740 => b:="6740";
                when 6741 => b:="6741";
                when 6742 => b:="6742";
                when 6743 => b:="6743";
                when 6744 => b:="6744";
                when 6745 => b:="6745";
                when 6746 => b:="6746";
                when 6747 => b:="6747";
                when 6748 => b:="6748";
                when 6749 => b:="6749";
                when 6750 => b:="6750";
                when 6751 => b:="6751";
                when 6752 => b:="6752";
                when 6753 => b:="6753";
                when 6754 => b:="6754";
                when 6755 => b:="6755";
                when 6756 => b:="6756";
                when 6757 => b:="6757";
                when 6758 => b:="6758";
                when 6759 => b:="6759";
                when 6760 => b:="6760";
                when 6761 => b:="6761";
                when 6762 => b:="6762";
                when 6763 => b:="6763";
                when 6764 => b:="6764";
                when 6765 => b:="6765";
                when 6766 => b:="6766";
                when 6767 => b:="6767";
                when 6768 => b:="6768";
                when 6769 => b:="6769";
                when 6770 => b:="6770";
                when 6771 => b:="6771";
                when 6772 => b:="6772";
                when 6773 => b:="6773";
                when 6774 => b:="6774";
                when 6775 => b:="6775";
                when 6776 => b:="6776";
                when 6777 => b:="6777";
                when 6778 => b:="6778";
                when 6779 => b:="6779";
                when 6780 => b:="6780";
                when 6781 => b:="6781";
                when 6782 => b:="6782";
                when 6783 => b:="6783";
                when 6784 => b:="6784";
                when 6785 => b:="6785";
                when 6786 => b:="6786";
                when 6787 => b:="6787";
                when 6788 => b:="6788";
                when 6789 => b:="6789";
                when 6790 => b:="6790";
                when 6791 => b:="6791";
                when 6792 => b:="6792";
                when 6793 => b:="6793";
                when 6794 => b:="6794";
                when 6795 => b:="6795";
                when 6796 => b:="6796";
                when 6797 => b:="6797";
                when 6798 => b:="6798";
                when 6799 => b:="6799";
                when 6800 => b:="6800";
                when 6801 => b:="6801";
                when 6802 => b:="6802";
                when 6803 => b:="6803";
                when 6804 => b:="6804";
                when 6805 => b:="6805";
                when 6806 => b:="6806";
                when 6807 => b:="6807";
                when 6808 => b:="6808";
                when 6809 => b:="6809";
                when 6810 => b:="6810";
                when 6811 => b:="6811";
                when 6812 => b:="6812";
                when 6813 => b:="6813";
                when 6814 => b:="6814";
                when 6815 => b:="6815";
                when 6816 => b:="6816";
                when 6817 => b:="6817";
                when 6818 => b:="6818";
                when 6819 => b:="6819";
                when 6820 => b:="6820";
                when 6821 => b:="6821";
                when 6822 => b:="6822";
                when 6823 => b:="6823";
                when 6824 => b:="6824";
                when 6825 => b:="6825";
                when 6826 => b:="6826";
                when 6827 => b:="6827";
                when 6828 => b:="6828";
                when 6829 => b:="6829";
                when 6830 => b:="6830";
                when 6831 => b:="6831";
                when 6832 => b:="6832";
                when 6833 => b:="6833";
                when 6834 => b:="6834";
                when 6835 => b:="6835";
                when 6836 => b:="6836";
                when 6837 => b:="6837";
                when 6838 => b:="6838";
                when 6839 => b:="6839";
                when 6840 => b:="6840";
                when 6841 => b:="6841";
                when 6842 => b:="6842";
                when 6843 => b:="6843";
                when 6844 => b:="6844";
                when 6845 => b:="6845";
                when 6846 => b:="6846";
                when 6847 => b:="6847";
                when 6848 => b:="6848";
                when 6849 => b:="6849";
                when 6850 => b:="6850";
                when 6851 => b:="6851";
                when 6852 => b:="6852";
                when 6853 => b:="6853";
                when 6854 => b:="6854";
                when 6855 => b:="6855";
                when 6856 => b:="6856";
                when 6857 => b:="6857";
                when 6858 => b:="6858";
                when 6859 => b:="6859";
                when 6860 => b:="6860";
                when 6861 => b:="6861";
                when 6862 => b:="6862";
                when 6863 => b:="6863";
                when 6864 => b:="6864";
                when 6865 => b:="6865";
                when 6866 => b:="6866";
                when 6867 => b:="6867";
                when 6868 => b:="6868";
                when 6869 => b:="6869";
                when 6870 => b:="6870";
                when 6871 => b:="6871";
                when 6872 => b:="6872";
                when 6873 => b:="6873";
                when 6874 => b:="6874";
                when 6875 => b:="6875";
                when 6876 => b:="6876";
                when 6877 => b:="6877";
                when 6878 => b:="6878";
                when 6879 => b:="6879";
                when 6880 => b:="6880";
                when 6881 => b:="6881";
                when 6882 => b:="6882";
                when 6883 => b:="6883";
                when 6884 => b:="6884";
                when 6885 => b:="6885";
                when 6886 => b:="6886";
                when 6887 => b:="6887";
                when 6888 => b:="6888";
                when 6889 => b:="6889";
                when 6890 => b:="6890";
                when 6891 => b:="6891";
                when 6892 => b:="6892";
                when 6893 => b:="6893";
                when 6894 => b:="6894";
                when 6895 => b:="6895";
                when 6896 => b:="6896";
                when 6897 => b:="6897";
                when 6898 => b:="6898";
                when 6899 => b:="6899";
                when 6900 => b:="6900";
                when 6901 => b:="6901";
                when 6902 => b:="6902";
                when 6903 => b:="6903";
                when 6904 => b:="6904";
                when 6905 => b:="6905";
                when 6906 => b:="6906";
                when 6907 => b:="6907";
                when 6908 => b:="6908";
                when 6909 => b:="6909";
                when 6910 => b:="6910";
                when 6911 => b:="6911";
                when 6912 => b:="6912";
                when 6913 => b:="6913";
                when 6914 => b:="6914";
                when 6915 => b:="6915";
                when 6916 => b:="6916";
                when 6917 => b:="6917";
                when 6918 => b:="6918";
                when 6919 => b:="6919";
                when 6920 => b:="6920";
                when 6921 => b:="6921";
                when 6922 => b:="6922";
                when 6923 => b:="6923";
                when 6924 => b:="6924";
                when 6925 => b:="6925";
                when 6926 => b:="6926";
                when 6927 => b:="6927";
                when 6928 => b:="6928";
                when 6929 => b:="6929";
                when 6930 => b:="6930";
                when 6931 => b:="6931";
                when 6932 => b:="6932";
                when 6933 => b:="6933";
                when 6934 => b:="6934";
                when 6935 => b:="6935";
                when 6936 => b:="6936";
                when 6937 => b:="6937";
                when 6938 => b:="6938";
                when 6939 => b:="6939";
                when 6940 => b:="6940";
                when 6941 => b:="6941";
                when 6942 => b:="6942";
                when 6943 => b:="6943";
                when 6944 => b:="6944";
                when 6945 => b:="6945";
                when 6946 => b:="6946";
                when 6947 => b:="6947";
                when 6948 => b:="6948";
                when 6949 => b:="6949";
                when 6950 => b:="6950";
                when 6951 => b:="6951";
                when 6952 => b:="6952";
                when 6953 => b:="6953";
                when 6954 => b:="6954";
                when 6955 => b:="6955";
                when 6956 => b:="6956";
                when 6957 => b:="6957";
                when 6958 => b:="6958";
                when 6959 => b:="6959";
                when 6960 => b:="6960";
                when 6961 => b:="6961";
                when 6962 => b:="6962";
                when 6963 => b:="6963";
                when 6964 => b:="6964";
                when 6965 => b:="6965";
                when 6966 => b:="6966";
                when 6967 => b:="6967";
                when 6968 => b:="6968";
                when 6969 => b:="6969";
                when 6970 => b:="6970";
                when 6971 => b:="6971";
                when 6972 => b:="6972";
                when 6973 => b:="6973";
                when 6974 => b:="6974";
                when 6975 => b:="6975";
                when 6976 => b:="6976";
                when 6977 => b:="6977";
                when 6978 => b:="6978";
                when 6979 => b:="6979";
                when 6980 => b:="6980";
                when 6981 => b:="6981";
                when 6982 => b:="6982";
                when 6983 => b:="6983";
                when 6984 => b:="6984";
                when 6985 => b:="6985";
                when 6986 => b:="6986";
                when 6987 => b:="6987";
                when 6988 => b:="6988";
                when 6989 => b:="6989";
                when 6990 => b:="6990";
                when 6991 => b:="6991";
                when 6992 => b:="6992";
                when 6993 => b:="6993";
                when 6994 => b:="6994";
                when 6995 => b:="6995";
                when 6996 => b:="6996";
                when 6997 => b:="6997";
                when 6998 => b:="6998";
                when 7000 => b:="7000";
                when 7001 => b:="7001";
                when 7002 => b:="7002";
                when 7003 => b:="7003";
                when 7004 => b:="7004";
                when 7005 => b:="7005";
                when 7006 => b:="7006";
                when 7007 => b:="7007";
                when 7008 => b:="7008";
                when 7009 => b:="7009";
                when 7010 => b:="7010";
                when 7011 => b:="7011";
                when 7012 => b:="7012";
                when 7013 => b:="7013";
                when 7014 => b:="7014";
                when 7015 => b:="7015";
                when 7016 => b:="7016";
                when 7017 => b:="7017";
                when 7018 => b:="7018";
                when 7019 => b:="7019";
                when 7020 => b:="7020";
                when 7021 => b:="7021";
                when 7022 => b:="7022";
                when 7023 => b:="7023";
                when 7024 => b:="7024";
                when 7025 => b:="7025";
                when 7026 => b:="7026";
                when 7027 => b:="7027";
                when 7028 => b:="7028";
                when 7029 => b:="7029";
                when 7030 => b:="7030";
                when 7031 => b:="7031";
                when 7032 => b:="7032";
                when 7033 => b:="7033";
                when 7034 => b:="7034";
                when 7035 => b:="7035";
                when 7036 => b:="7036";
                when 7037 => b:="7037";
                when 7038 => b:="7038";
                when 7039 => b:="7039";
                when 7040 => b:="7040";
                when 7041 => b:="7041";
                when 7042 => b:="7042";
                when 7043 => b:="7043";
                when 7044 => b:="7044";
                when 7045 => b:="7045";
                when 7046 => b:="7046";
                when 7047 => b:="7047";
                when 7048 => b:="7048";
                when 7049 => b:="7049";
                when 7050 => b:="7050";
                when 7051 => b:="7051";
                when 7052 => b:="7052";
                when 7053 => b:="7053";
                when 7054 => b:="7054";
                when 7055 => b:="7055";
                when 7056 => b:="7056";
                when 7057 => b:="7057";
                when 7058 => b:="7058";
                when 7059 => b:="7059";
                when 7060 => b:="7060";
                when 7061 => b:="7061";
                when 7062 => b:="7062";
                when 7063 => b:="7063";
                when 7064 => b:="7064";
                when 7065 => b:="7065";
                when 7066 => b:="7066";
                when 7067 => b:="7067";
                when 7068 => b:="7068";
                when 7069 => b:="7069";
                when 7070 => b:="7070";
                when 7071 => b:="7071";
                when 7072 => b:="7072";
                when 7073 => b:="7073";
                when 7074 => b:="7074";
                when 7075 => b:="7075";
                when 7076 => b:="7076";
                when 7077 => b:="7077";
                when 7078 => b:="7078";
                when 7079 => b:="7079";
                when 7080 => b:="7080";
                when 7081 => b:="7081";
                when 7082 => b:="7082";
                when 7083 => b:="7083";
                when 7084 => b:="7084";
                when 7085 => b:="7085";
                when 7086 => b:="7086";
                when 7087 => b:="7087";
                when 7088 => b:="7088";
                when 7089 => b:="7089";
                when 7090 => b:="7090";
                when 7091 => b:="7091";
                when 7092 => b:="7092";
                when 7093 => b:="7093";
                when 7094 => b:="7094";
                when 7095 => b:="7095";
                when 7096 => b:="7096";
                when 7097 => b:="7097";
                when 7098 => b:="7098";
                when 7099 => b:="7099";
                when 7100 => b:="7100";
                when 7101 => b:="7101";
                when 7102 => b:="7102";
                when 7103 => b:="7103";
                when 7104 => b:="7104";
                when 7105 => b:="7105";
                when 7106 => b:="7106";
                when 7107 => b:="7107";
                when 7108 => b:="7108";
                when 7109 => b:="7109";
                when 7110 => b:="7110";
                when 7111 => b:="7111";
                when 7112 => b:="7112";
                when 7113 => b:="7113";
                when 7114 => b:="7114";
                when 7115 => b:="7115";
                when 7116 => b:="7116";
                when 7117 => b:="7117";
                when 7118 => b:="7118";
                when 7119 => b:="7119";
                when 7120 => b:="7120";
                when 7121 => b:="7121";
                when 7122 => b:="7122";
                when 7123 => b:="7123";
                when 7124 => b:="7124";
                when 7125 => b:="7125";
                when 7126 => b:="7126";
                when 7127 => b:="7127";
                when 7128 => b:="7128";
                when 7129 => b:="7129";
                when 7130 => b:="7130";
                when 7131 => b:="7131";
                when 7132 => b:="7132";
                when 7133 => b:="7133";
                when 7134 => b:="7134";
                when 7135 => b:="7135";
                when 7136 => b:="7136";
                when 7137 => b:="7137";
                when 7138 => b:="7138";
                when 7139 => b:="7139";
                when 7140 => b:="7140";
                when 7141 => b:="7141";
                when 7142 => b:="7142";
                when 7143 => b:="7143";
                when 7144 => b:="7144";
                when 7145 => b:="7145";
                when 7146 => b:="7146";
                when 7147 => b:="7147";
                when 7148 => b:="7148";
                when 7149 => b:="7149";
                when 7150 => b:="7150";
                when 7151 => b:="7151";
                when 7152 => b:="7152";
                when 7153 => b:="7153";
                when 7154 => b:="7154";
                when 7155 => b:="7155";
                when 7156 => b:="7156";
                when 7157 => b:="7157";
                when 7158 => b:="7158";
                when 7159 => b:="7159";
                when 7160 => b:="7160";
                when 7161 => b:="7161";
                when 7162 => b:="7162";
                when 7163 => b:="7163";
                when 7164 => b:="7164";
                when 7165 => b:="7165";
                when 7166 => b:="7166";
                when 7167 => b:="7167";
                when 7168 => b:="7168";
                when 7169 => b:="7169";
                when 7170 => b:="7170";
                when 7171 => b:="7171";
                when 7172 => b:="7172";
                when 7173 => b:="7173";
                when 7174 => b:="7174";
                when 7175 => b:="7175";
                when 7176 => b:="7176";
                when 7177 => b:="7177";
                when 7178 => b:="7178";
                when 7179 => b:="7179";
                when 7180 => b:="7180";
                when 7181 => b:="7181";
                when 7182 => b:="7182";
                when 7183 => b:="7183";
                when 7184 => b:="7184";
                when 7185 => b:="7185";
                when 7186 => b:="7186";
                when 7187 => b:="7187";
                when 7188 => b:="7188";
                when 7189 => b:="7189";
                when 7190 => b:="7190";
                when 7191 => b:="7191";
                when 7192 => b:="7192";
                when 7193 => b:="7193";
                when 7194 => b:="7194";
                when 7195 => b:="7195";
                when 7196 => b:="7196";
                when 7197 => b:="7197";
                when 7198 => b:="7198";
                when 7199 => b:="7199";
                when 7200 => b:="7200";
                when 7201 => b:="7201";
                when 7202 => b:="7202";
                when 7203 => b:="7203";
                when 7204 => b:="7204";
                when 7205 => b:="7205";
                when 7206 => b:="7206";
                when 7207 => b:="7207";
                when 7208 => b:="7208";
                when 7209 => b:="7209";
                when 7210 => b:="7210";
                when 7211 => b:="7211";
                when 7212 => b:="7212";
                when 7213 => b:="7213";
                when 7214 => b:="7214";
                when 7215 => b:="7215";
                when 7216 => b:="7216";
                when 7217 => b:="7217";
                when 7218 => b:="7218";
                when 7219 => b:="7219";
                when 7220 => b:="7220";
                when 7221 => b:="7221";
                when 7222 => b:="7222";
                when 7223 => b:="7223";
                when 7224 => b:="7224";
                when 7225 => b:="7225";
                when 7226 => b:="7226";
                when 7227 => b:="7227";
                when 7228 => b:="7228";
                when 7229 => b:="7229";
                when 7230 => b:="7230";
                when 7231 => b:="7231";
                when 7232 => b:="7232";
                when 7233 => b:="7233";
                when 7234 => b:="7234";
                when 7235 => b:="7235";
                when 7236 => b:="7236";
                when 7237 => b:="7237";
                when 7238 => b:="7238";
                when 7239 => b:="7239";
                when 7240 => b:="7240";
                when 7241 => b:="7241";
                when 7242 => b:="7242";
                when 7243 => b:="7243";
                when 7244 => b:="7244";
                when 7245 => b:="7245";
                when 7246 => b:="7246";
                when 7247 => b:="7247";
                when 7248 => b:="7248";
                when 7249 => b:="7249";
                when 7250 => b:="7250";
                when 7251 => b:="7251";
                when 7252 => b:="7252";
                when 7253 => b:="7253";
                when 7254 => b:="7254";
                when 7255 => b:="7255";
                when 7256 => b:="7256";
                when 7257 => b:="7257";
                when 7258 => b:="7258";
                when 7259 => b:="7259";
                when 7260 => b:="7260";
                when 7261 => b:="7261";
                when 7262 => b:="7262";
                when 7263 => b:="7263";
                when 7264 => b:="7264";
                when 7265 => b:="7265";
                when 7266 => b:="7266";
                when 7267 => b:="7267";
                when 7268 => b:="7268";
                when 7269 => b:="7269";
                when 7270 => b:="7270";
                when 7271 => b:="7271";
                when 7272 => b:="7272";
                when 7273 => b:="7273";
                when 7274 => b:="7274";
                when 7275 => b:="7275";
                when 7276 => b:="7276";
                when 7277 => b:="7277";
                when 7278 => b:="7278";
                when 7279 => b:="7279";
                when 7280 => b:="7280";
                when 7281 => b:="7281";
                when 7282 => b:="7282";
                when 7283 => b:="7283";
                when 7284 => b:="7284";
                when 7285 => b:="7285";
                when 7286 => b:="7286";
                when 7287 => b:="7287";
                when 7288 => b:="7288";
                when 7289 => b:="7289";
                when 7290 => b:="7290";
                when 7291 => b:="7291";
                when 7292 => b:="7292";
                when 7293 => b:="7293";
                when 7294 => b:="7294";
                when 7295 => b:="7295";
                when 7296 => b:="7296";
                when 7297 => b:="7297";
                when 7298 => b:="7298";
                when 7299 => b:="7299";
                when 7300 => b:="7300";
                when 7301 => b:="7301";
                when 7302 => b:="7302";
                when 7303 => b:="7303";
                when 7304 => b:="7304";
                when 7305 => b:="7305";
                when 7306 => b:="7306";
                when 7307 => b:="7307";
                when 7308 => b:="7308";
                when 7309 => b:="7309";
                when 7310 => b:="7310";
                when 7311 => b:="7311";
                when 7312 => b:="7312";
                when 7313 => b:="7313";
                when 7314 => b:="7314";
                when 7315 => b:="7315";
                when 7316 => b:="7316";
                when 7317 => b:="7317";
                when 7318 => b:="7318";
                when 7319 => b:="7319";
                when 7320 => b:="7320";
                when 7321 => b:="7321";
                when 7322 => b:="7322";
                when 7323 => b:="7323";
                when 7324 => b:="7324";
                when 7325 => b:="7325";
                when 7326 => b:="7326";
                when 7327 => b:="7327";
                when 7328 => b:="7328";
                when 7329 => b:="7329";
                when 7330 => b:="7330";
                when 7331 => b:="7331";
                when 7332 => b:="7332";
                when 7333 => b:="7333";
                when 7334 => b:="7334";
                when 7335 => b:="7335";
                when 7336 => b:="7336";
                when 7337 => b:="7337";
                when 7338 => b:="7338";
                when 7339 => b:="7339";
                when 7340 => b:="7340";
                when 7341 => b:="7341";
                when 7342 => b:="7342";
                when 7343 => b:="7343";
                when 7344 => b:="7344";
                when 7345 => b:="7345";
                when 7346 => b:="7346";
                when 7347 => b:="7347";
                when 7348 => b:="7348";
                when 7349 => b:="7349";
                when 7350 => b:="7350";
                when 7351 => b:="7351";
                when 7352 => b:="7352";
                when 7353 => b:="7353";
                when 7354 => b:="7354";
                when 7355 => b:="7355";
                when 7356 => b:="7356";
                when 7357 => b:="7357";
                when 7358 => b:="7358";
                when 7359 => b:="7359";
                when 7360 => b:="7360";
                when 7361 => b:="7361";
                when 7362 => b:="7362";
                when 7363 => b:="7363";
                when 7364 => b:="7364";
                when 7365 => b:="7365";
                when 7366 => b:="7366";
                when 7367 => b:="7367";
                when 7368 => b:="7368";
                when 7369 => b:="7369";
                when 7370 => b:="7370";
                when 7371 => b:="7371";
                when 7372 => b:="7372";
                when 7373 => b:="7373";
                when 7374 => b:="7374";
                when 7375 => b:="7375";
                when 7376 => b:="7376";
                when 7377 => b:="7377";
                when 7378 => b:="7378";
                when 7379 => b:="7379";
                when 7380 => b:="7380";
                when 7381 => b:="7381";
                when 7382 => b:="7382";
                when 7383 => b:="7383";
                when 7384 => b:="7384";
                when 7385 => b:="7385";
                when 7386 => b:="7386";
                when 7387 => b:="7387";
                when 7388 => b:="7388";
                when 7389 => b:="7389";
                when 7390 => b:="7390";
                when 7391 => b:="7391";
                when 7392 => b:="7392";
                when 7393 => b:="7393";
                when 7394 => b:="7394";
                when 7395 => b:="7395";
                when 7396 => b:="7396";
                when 7397 => b:="7397";
                when 7398 => b:="7398";
                when 7399 => b:="7399";
                when 7400 => b:="7400";
                when 7401 => b:="7401";
                when 7402 => b:="7402";
                when 7403 => b:="7403";
                when 7404 => b:="7404";
                when 7405 => b:="7405";
                when 7406 => b:="7406";
                when 7407 => b:="7407";
                when 7408 => b:="7408";
                when 7409 => b:="7409";
                when 7410 => b:="7410";
                when 7411 => b:="7411";
                when 7412 => b:="7412";
                when 7413 => b:="7413";
                when 7414 => b:="7414";
                when 7415 => b:="7415";
                when 7416 => b:="7416";
                when 7417 => b:="7417";
                when 7418 => b:="7418";
                when 7419 => b:="7419";
                when 7420 => b:="7420";
                when 7421 => b:="7421";
                when 7422 => b:="7422";
                when 7423 => b:="7423";
                when 7424 => b:="7424";
                when 7425 => b:="7425";
                when 7426 => b:="7426";
                when 7427 => b:="7427";
                when 7428 => b:="7428";
                when 7429 => b:="7429";
                when 7430 => b:="7430";
                when 7431 => b:="7431";
                when 7432 => b:="7432";
                when 7433 => b:="7433";
                when 7434 => b:="7434";
                when 7435 => b:="7435";
                when 7436 => b:="7436";
                when 7437 => b:="7437";
                when 7438 => b:="7438";
                when 7439 => b:="7439";
                when 7440 => b:="7440";
                when 7441 => b:="7441";
                when 7442 => b:="7442";
                when 7443 => b:="7443";
                when 7444 => b:="7444";
                when 7445 => b:="7445";
                when 7446 => b:="7446";
                when 7447 => b:="7447";
                when 7448 => b:="7448";
                when 7449 => b:="7449";
                when 7450 => b:="7450";
                when 7451 => b:="7451";
                when 7452 => b:="7452";
                when 7453 => b:="7453";
                when 7454 => b:="7454";
                when 7455 => b:="7455";
                when 7456 => b:="7456";
                when 7457 => b:="7457";
                when 7458 => b:="7458";
                when 7459 => b:="7459";
                when 7460 => b:="7460";
                when 7461 => b:="7461";
                when 7462 => b:="7462";
                when 7463 => b:="7463";
                when 7464 => b:="7464";
                when 7465 => b:="7465";
                when 7466 => b:="7466";
                when 7467 => b:="7467";
                when 7468 => b:="7468";
                when 7469 => b:="7469";
                when 7470 => b:="7470";
                when 7471 => b:="7471";
                when 7472 => b:="7472";
                when 7473 => b:="7473";
                when 7474 => b:="7474";
                when 7475 => b:="7475";
                when 7476 => b:="7476";
                when 7477 => b:="7477";
                when 7478 => b:="7478";
                when 7479 => b:="7479";
                when 7480 => b:="7480";
                when 7481 => b:="7481";
                when 7482 => b:="7482";
                when 7483 => b:="7483";
                when 7484 => b:="7484";
                when 7485 => b:="7485";
                when 7486 => b:="7486";
                when 7487 => b:="7487";
                when 7488 => b:="7488";
                when 7489 => b:="7489";
                when 7490 => b:="7490";
                when 7491 => b:="7491";
                when 7492 => b:="7492";
                when 7493 => b:="7493";
                when 7494 => b:="7494";
                when 7495 => b:="7495";
                when 7496 => b:="7496";
                when 7497 => b:="7497";
                when 7498 => b:="7498";
                when 7499 => b:="7499";
                when 7500 => b:="7500";
                when 7501 => b:="7501";
                when 7502 => b:="7502";
                when 7503 => b:="7503";
                when 7504 => b:="7504";
                when 7505 => b:="7505";
                when 7506 => b:="7506";
                when 7507 => b:="7507";
                when 7508 => b:="7508";
                when 7509 => b:="7509";
                when 7510 => b:="7510";
                when 7511 => b:="7511";
                when 7512 => b:="7512";
                when 7513 => b:="7513";
                when 7514 => b:="7514";
                when 7515 => b:="7515";
                when 7516 => b:="7516";
                when 7517 => b:="7517";
                when 7518 => b:="7518";
                when 7519 => b:="7519";
                when 7520 => b:="7520";
                when 7521 => b:="7521";
                when 7522 => b:="7522";
                when 7523 => b:="7523";
                when 7524 => b:="7524";
                when 7525 => b:="7525";
                when 7526 => b:="7526";
                when 7527 => b:="7527";
                when 7528 => b:="7528";
                when 7529 => b:="7529";
                when 7530 => b:="7530";
                when 7531 => b:="7531";
                when 7532 => b:="7532";
                when 7533 => b:="7533";
                when 7534 => b:="7534";
                when 7535 => b:="7535";
                when 7536 => b:="7536";
                when 7537 => b:="7537";
                when 7538 => b:="7538";
                when 7539 => b:="7539";
                when 7540 => b:="7540";
                when 7541 => b:="7541";
                when 7542 => b:="7542";
                when 7543 => b:="7543";
                when 7544 => b:="7544";
                when 7545 => b:="7545";
                when 7546 => b:="7546";
                when 7547 => b:="7547";
                when 7548 => b:="7548";
                when 7549 => b:="7549";
                when 7550 => b:="7550";
                when 7551 => b:="7551";
                when 7552 => b:="7552";
                when 7553 => b:="7553";
                when 7554 => b:="7554";
                when 7555 => b:="7555";
                when 7556 => b:="7556";
                when 7557 => b:="7557";
                when 7558 => b:="7558";
                when 7559 => b:="7559";
                when 7560 => b:="7560";
                when 7561 => b:="7561";
                when 7562 => b:="7562";
                when 7563 => b:="7563";
                when 7564 => b:="7564";
                when 7565 => b:="7565";
                when 7566 => b:="7566";
                when 7567 => b:="7567";
                when 7568 => b:="7568";
                when 7569 => b:="7569";
                when 7570 => b:="7570";
                when 7571 => b:="7571";
                when 7572 => b:="7572";
                when 7573 => b:="7573";
                when 7574 => b:="7574";
                when 7575 => b:="7575";
                when 7576 => b:="7576";
                when 7577 => b:="7577";
                when 7578 => b:="7578";
                when 7579 => b:="7579";
                when 7580 => b:="7580";
                when 7581 => b:="7581";
                when 7582 => b:="7582";
                when 7583 => b:="7583";
                when 7584 => b:="7584";
                when 7585 => b:="7585";
                when 7586 => b:="7586";
                when 7587 => b:="7587";
                when 7588 => b:="7588";
                when 7589 => b:="7589";
                when 7590 => b:="7590";
                when 7591 => b:="7591";
                when 7592 => b:="7592";
                when 7593 => b:="7593";
                when 7594 => b:="7594";
                when 7595 => b:="7595";
                when 7596 => b:="7596";
                when 7597 => b:="7597";
                when 7598 => b:="7598";
                when 7599 => b:="7599";
                when 7600 => b:="7600";
                when 7601 => b:="7601";
                when 7602 => b:="7602";
                when 7603 => b:="7603";
                when 7604 => b:="7604";
                when 7605 => b:="7605";
                when 7606 => b:="7606";
                when 7607 => b:="7607";
                when 7608 => b:="7608";
                when 7609 => b:="7609";
                when 7610 => b:="7610";
                when 7611 => b:="7611";
                when 7612 => b:="7612";
                when 7613 => b:="7613";
                when 7614 => b:="7614";
                when 7615 => b:="7615";
                when 7616 => b:="7616";
                when 7617 => b:="7617";
                when 7618 => b:="7618";
                when 7619 => b:="7619";
                when 7620 => b:="7620";
                when 7621 => b:="7621";
                when 7622 => b:="7622";
                when 7623 => b:="7623";
                when 7624 => b:="7624";
                when 7625 => b:="7625";
                when 7626 => b:="7626";
                when 7627 => b:="7627";
                when 7628 => b:="7628";
                when 7629 => b:="7629";
                when 7630 => b:="7630";
                when 7631 => b:="7631";
                when 7632 => b:="7632";
                when 7633 => b:="7633";
                when 7634 => b:="7634";
                when 7635 => b:="7635";
                when 7636 => b:="7636";
                when 7637 => b:="7637";
                when 7638 => b:="7638";
                when 7639 => b:="7639";
                when 7640 => b:="7640";
                when 7641 => b:="7641";
                when 7642 => b:="7642";
                when 7643 => b:="7643";
                when 7644 => b:="7644";
                when 7645 => b:="7645";
                when 7646 => b:="7646";
                when 7647 => b:="7647";
                when 7648 => b:="7648";
                when 7649 => b:="7649";
                when 7650 => b:="7650";
                when 7651 => b:="7651";
                when 7652 => b:="7652";
                when 7653 => b:="7653";
                when 7654 => b:="7654";
                when 7655 => b:="7655";
                when 7656 => b:="7656";
                when 7657 => b:="7657";
                when 7658 => b:="7658";
                when 7659 => b:="7659";
                when 7660 => b:="7660";
                when 7661 => b:="7661";
                when 7662 => b:="7662";
                when 7663 => b:="7663";
                when 7664 => b:="7664";
                when 7665 => b:="7665";
                when 7666 => b:="7666";
                when 7667 => b:="7667";
                when 7668 => b:="7668";
                when 7669 => b:="7669";
                when 7670 => b:="7670";
                when 7671 => b:="7671";
                when 7672 => b:="7672";
                when 7673 => b:="7673";
                when 7674 => b:="7674";
                when 7675 => b:="7675";
                when 7676 => b:="7676";
                when 7677 => b:="7677";
                when 7678 => b:="7678";
                when 7679 => b:="7679";
                when 7680 => b:="7680";
                when 7681 => b:="7681";
                when 7682 => b:="7682";
                when 7683 => b:="7683";
                when 7684 => b:="7684";
                when 7685 => b:="7685";
                when 7686 => b:="7686";
                when 7687 => b:="7687";
                when 7688 => b:="7688";
                when 7689 => b:="7689";
                when 7690 => b:="7690";
                when 7691 => b:="7691";
                when 7692 => b:="7692";
                when 7693 => b:="7693";
                when 7694 => b:="7694";
                when 7695 => b:="7695";
                when 7696 => b:="7696";
                when 7697 => b:="7697";
                when 7698 => b:="7698";
                when 7699 => b:="7699";
                when 7700 => b:="7700";
                when 7701 => b:="7701";
                when 7702 => b:="7702";
                when 7703 => b:="7703";
                when 7704 => b:="7704";
                when 7705 => b:="7705";
                when 7706 => b:="7706";
                when 7707 => b:="7707";
                when 7708 => b:="7708";
                when 7709 => b:="7709";
                when 7710 => b:="7710";
                when 7711 => b:="7711";
                when 7712 => b:="7712";
                when 7713 => b:="7713";
                when 7714 => b:="7714";
                when 7715 => b:="7715";
                when 7716 => b:="7716";
                when 7717 => b:="7717";
                when 7718 => b:="7718";
                when 7719 => b:="7719";
                when 7720 => b:="7720";
                when 7721 => b:="7721";
                when 7722 => b:="7722";
                when 7723 => b:="7723";
                when 7724 => b:="7724";
                when 7725 => b:="7725";
                when 7726 => b:="7726";
                when 7727 => b:="7727";
                when 7728 => b:="7728";
                when 7729 => b:="7729";
                when 7730 => b:="7730";
                when 7731 => b:="7731";
                when 7732 => b:="7732";
                when 7733 => b:="7733";
                when 7734 => b:="7734";
                when 7735 => b:="7735";
                when 7736 => b:="7736";
                when 7737 => b:="7737";
                when 7738 => b:="7738";
                when 7739 => b:="7739";
                when 7740 => b:="7740";
                when 7741 => b:="7741";
                when 7742 => b:="7742";
                when 7743 => b:="7743";
                when 7744 => b:="7744";
                when 7745 => b:="7745";
                when 7746 => b:="7746";
                when 7747 => b:="7747";
                when 7748 => b:="7748";
                when 7749 => b:="7749";
                when 7750 => b:="7750";
                when 7751 => b:="7751";
                when 7752 => b:="7752";
                when 7753 => b:="7753";
                when 7754 => b:="7754";
                when 7755 => b:="7755";
                when 7756 => b:="7756";
                when 7757 => b:="7757";
                when 7758 => b:="7758";
                when 7759 => b:="7759";
                when 7760 => b:="7760";
                when 7761 => b:="7761";
                when 7762 => b:="7762";
                when 7763 => b:="7763";
                when 7764 => b:="7764";
                when 7765 => b:="7765";
                when 7766 => b:="7766";
                when 7767 => b:="7767";
                when 7768 => b:="7768";
                when 7769 => b:="7769";
                when 7770 => b:="7770";
                when 7771 => b:="7771";
                when 7772 => b:="7772";
                when 7773 => b:="7773";
                when 7774 => b:="7774";
                when 7775 => b:="7775";
                when 7776 => b:="7776";
                when 7777 => b:="7777";
                when 7778 => b:="7778";
                when 7779 => b:="7779";
                when 7780 => b:="7780";
                when 7781 => b:="7781";
                when 7782 => b:="7782";
                when 7783 => b:="7783";
                when 7784 => b:="7784";
                when 7785 => b:="7785";
                when 7786 => b:="7786";
                when 7787 => b:="7787";
                when 7788 => b:="7788";
                when 7789 => b:="7789";
                when 7790 => b:="7790";
                when 7791 => b:="7791";
                when 7792 => b:="7792";
                when 7793 => b:="7793";
                when 7794 => b:="7794";
                when 7795 => b:="7795";
                when 7796 => b:="7796";
                when 7797 => b:="7797";
                when 7798 => b:="7798";
                when 7799 => b:="7799";
                when 7800 => b:="7800";
                when 7801 => b:="7801";
                when 7802 => b:="7802";
                when 7803 => b:="7803";
                when 7804 => b:="7804";
                when 7805 => b:="7805";
                when 7806 => b:="7806";
                when 7807 => b:="7807";
                when 7808 => b:="7808";
                when 7809 => b:="7809";
                when 7810 => b:="7810";
                when 7811 => b:="7811";
                when 7812 => b:="7812";
                when 7813 => b:="7813";
                when 7814 => b:="7814";
                when 7815 => b:="7815";
                when 7816 => b:="7816";
                when 7817 => b:="7817";
                when 7818 => b:="7818";
                when 7819 => b:="7819";
                when 7820 => b:="7820";
                when 7821 => b:="7821";
                when 7822 => b:="7822";
                when 7823 => b:="7823";
                when 7824 => b:="7824";
                when 7825 => b:="7825";
                when 7826 => b:="7826";
                when 7827 => b:="7827";
                when 7828 => b:="7828";
                when 7829 => b:="7829";
                when 7830 => b:="7830";
                when 7831 => b:="7831";
                when 7832 => b:="7832";
                when 7833 => b:="7833";
                when 7834 => b:="7834";
                when 7835 => b:="7835";
                when 7836 => b:="7836";
                when 7837 => b:="7837";
                when 7838 => b:="7838";
                when 7839 => b:="7839";
                when 7840 => b:="7840";
                when 7841 => b:="7841";
                when 7842 => b:="7842";
                when 7843 => b:="7843";
                when 7844 => b:="7844";
                when 7845 => b:="7845";
                when 7846 => b:="7846";
                when 7847 => b:="7847";
                when 7848 => b:="7848";
                when 7849 => b:="7849";
                when 7850 => b:="7850";
                when 7851 => b:="7851";
                when 7852 => b:="7852";
                when 7853 => b:="7853";
                when 7854 => b:="7854";
                when 7855 => b:="7855";
                when 7856 => b:="7856";
                when 7857 => b:="7857";
                when 7858 => b:="7858";
                when 7859 => b:="7859";
                when 7860 => b:="7860";
                when 7861 => b:="7861";
                when 7862 => b:="7862";
                when 7863 => b:="7863";
                when 7864 => b:="7864";
                when 7865 => b:="7865";
                when 7866 => b:="7866";
                when 7867 => b:="7867";
                when 7868 => b:="7868";
                when 7869 => b:="7869";
                when 7870 => b:="7870";
                when 7871 => b:="7871";
                when 7872 => b:="7872";
                when 7873 => b:="7873";
                when 7874 => b:="7874";
                when 7875 => b:="7875";
                when 7876 => b:="7876";
                when 7877 => b:="7877";
                when 7878 => b:="7878";
                when 7879 => b:="7879";
                when 7880 => b:="7880";
                when 7881 => b:="7881";
                when 7882 => b:="7882";
                when 7883 => b:="7883";
                when 7884 => b:="7884";
                when 7885 => b:="7885";
                when 7886 => b:="7886";
                when 7887 => b:="7887";
                when 7888 => b:="7888";
                when 7889 => b:="7889";
                when 7890 => b:="7890";
                when 7891 => b:="7891";
                when 7892 => b:="7892";
                when 7893 => b:="7893";
                when 7894 => b:="7894";
                when 7895 => b:="7895";
                when 7896 => b:="7896";
                when 7897 => b:="7897";
                when 7898 => b:="7898";
                when 7899 => b:="7899";
                when 7900 => b:="7900";
                when 7901 => b:="7901";
                when 7902 => b:="7902";
                when 7903 => b:="7903";
                when 7904 => b:="7904";
                when 7905 => b:="7905";
                when 7906 => b:="7906";
                when 7907 => b:="7907";
                when 7908 => b:="7908";
                when 7909 => b:="7909";
                when 7910 => b:="7910";
                when 7911 => b:="7911";
                when 7912 => b:="7912";
                when 7913 => b:="7913";
                when 7914 => b:="7914";
                when 7915 => b:="7915";
                when 7916 => b:="7916";
                when 7917 => b:="7917";
                when 7918 => b:="7918";
                when 7919 => b:="7919";
                when 7920 => b:="7920";
                when 7921 => b:="7921";
                when 7922 => b:="7922";
                when 7923 => b:="7923";
                when 7924 => b:="7924";
                when 7925 => b:="7925";
                when 7926 => b:="7926";
                when 7927 => b:="7927";
                when 7928 => b:="7928";
                when 7929 => b:="7929";
                when 7930 => b:="7930";
                when 7931 => b:="7931";
                when 7932 => b:="7932";
                when 7933 => b:="7933";
                when 7934 => b:="7934";
                when 7935 => b:="7935";
                when 7936 => b:="7936";
                when 7937 => b:="7937";
                when 7938 => b:="7938";
                when 7939 => b:="7939";
                when 7940 => b:="7940";
                when 7941 => b:="7941";
                when 7942 => b:="7942";
                when 7943 => b:="7943";
                when 7944 => b:="7944";
                when 7945 => b:="7945";
                when 7946 => b:="7946";
                when 7947 => b:="7947";
                when 7948 => b:="7948";
                when 7949 => b:="7949";
                when 7950 => b:="7950";
                when 7951 => b:="7951";
                when 7952 => b:="7952";
                when 7953 => b:="7953";
                when 7954 => b:="7954";
                when 7955 => b:="7955";
                when 7956 => b:="7956";
                when 7957 => b:="7957";
                when 7958 => b:="7958";
                when 7959 => b:="7959";
                when 7960 => b:="7960";
                when 7961 => b:="7961";
                when 7962 => b:="7962";
                when 7963 => b:="7963";
                when 7964 => b:="7964";
                when 7965 => b:="7965";
                when 7966 => b:="7966";
                when 7967 => b:="7967";
                when 7968 => b:="7968";
                when 7969 => b:="7969";
                when 7970 => b:="7970";
                when 7971 => b:="7971";
                when 7972 => b:="7972";
                when 7973 => b:="7973";
                when 7974 => b:="7974";
                when 7975 => b:="7975";
                when 7976 => b:="7976";
                when 7977 => b:="7977";
                when 7978 => b:="7978";
                when 7979 => b:="7979";
                when 7980 => b:="7980";
                when 7981 => b:="7981";
                when 7982 => b:="7982";
                when 7983 => b:="7983";
                when 7984 => b:="7984";
                when 7985 => b:="7985";
                when 7986 => b:="7986";
                when 7987 => b:="7987";
                when 7988 => b:="7988";
                when 7989 => b:="7989";
                when 7990 => b:="7990";
                when 7991 => b:="7991";
                when 7992 => b:="7992";
                when 7993 => b:="7993";
                when 7994 => b:="7994";
                when 7995 => b:="7995";
                when 7996 => b:="7996";
                when 7997 => b:="7997";
                when 7998 => b:="7998";
                when 8000 => b:="8000";
                when 8001 => b:="8001";
                when 8002 => b:="8002";
                when 8003 => b:="8003";
                when 8004 => b:="8004";
                when 8005 => b:="8005";
                when 8006 => b:="8006";
                when 8007 => b:="8007";
                when 8008 => b:="8008";
                when 8009 => b:="8009";
                when 8010 => b:="8010";
                when 8011 => b:="8011";
                when 8012 => b:="8012";
                when 8013 => b:="8013";
                when 8014 => b:="8014";
                when 8015 => b:="8015";
                when 8016 => b:="8016";
                when 8017 => b:="8017";
                when 8018 => b:="8018";
                when 8019 => b:="8019";
                when 8020 => b:="8020";
                when 8021 => b:="8021";
                when 8022 => b:="8022";
                when 8023 => b:="8023";
                when 8024 => b:="8024";
                when 8025 => b:="8025";
                when 8026 => b:="8026";
                when 8027 => b:="8027";
                when 8028 => b:="8028";
                when 8029 => b:="8029";
                when 8030 => b:="8030";
                when 8031 => b:="8031";
                when 8032 => b:="8032";
                when 8033 => b:="8033";
                when 8034 => b:="8034";
                when 8035 => b:="8035";
                when 8036 => b:="8036";
                when 8037 => b:="8037";
                when 8038 => b:="8038";
                when 8039 => b:="8039";
                when 8040 => b:="8040";
                when 8041 => b:="8041";
                when 8042 => b:="8042";
                when 8043 => b:="8043";
                when 8044 => b:="8044";
                when 8045 => b:="8045";
                when 8046 => b:="8046";
                when 8047 => b:="8047";
                when 8048 => b:="8048";
                when 8049 => b:="8049";
                when 8050 => b:="8050";
                when 8051 => b:="8051";
                when 8052 => b:="8052";
                when 8053 => b:="8053";
                when 8054 => b:="8054";
                when 8055 => b:="8055";
                when 8056 => b:="8056";
                when 8057 => b:="8057";
                when 8058 => b:="8058";
                when 8059 => b:="8059";
                when 8060 => b:="8060";
                when 8061 => b:="8061";
                when 8062 => b:="8062";
                when 8063 => b:="8063";
                when 8064 => b:="8064";
                when 8065 => b:="8065";
                when 8066 => b:="8066";
                when 8067 => b:="8067";
                when 8068 => b:="8068";
                when 8069 => b:="8069";
                when 8070 => b:="8070";
                when 8071 => b:="8071";
                when 8072 => b:="8072";
                when 8073 => b:="8073";
                when 8074 => b:="8074";
                when 8075 => b:="8075";
                when 8076 => b:="8076";
                when 8077 => b:="8077";
                when 8078 => b:="8078";
                when 8079 => b:="8079";
                when 8080 => b:="8080";
                when 8081 => b:="8081";
                when 8082 => b:="8082";
                when 8083 => b:="8083";
                when 8084 => b:="8084";
                when 8085 => b:="8085";
                when 8086 => b:="8086";
                when 8087 => b:="8087";
                when 8088 => b:="8088";
                when 8089 => b:="8089";
                when 8090 => b:="8090";
                when 8091 => b:="8091";
                when 8092 => b:="8092";
                when 8093 => b:="8093";
                when 8094 => b:="8094";
                when 8095 => b:="8095";
                when 8096 => b:="8096";
                when 8097 => b:="8097";
                when 8098 => b:="8098";
                when 8099 => b:="8099";
                when 8100 => b:="8100";
                when 8101 => b:="8101";
                when 8102 => b:="8102";
                when 8103 => b:="8103";
                when 8104 => b:="8104";
                when 8105 => b:="8105";
                when 8106 => b:="8106";
                when 8107 => b:="8107";
                when 8108 => b:="8108";
                when 8109 => b:="8109";
                when 8110 => b:="8110";
                when 8111 => b:="8111";
                when 8112 => b:="8112";
                when 8113 => b:="8113";
                when 8114 => b:="8114";
                when 8115 => b:="8115";
                when 8116 => b:="8116";
                when 8117 => b:="8117";
                when 8118 => b:="8118";
                when 8119 => b:="8119";
                when 8120 => b:="8120";
                when 8121 => b:="8121";
                when 8122 => b:="8122";
                when 8123 => b:="8123";
                when 8124 => b:="8124";
                when 8125 => b:="8125";
                when 8126 => b:="8126";
                when 8127 => b:="8127";
                when 8128 => b:="8128";
                when 8129 => b:="8129";
                when 8130 => b:="8130";
                when 8131 => b:="8131";
                when 8132 => b:="8132";
                when 8133 => b:="8133";
                when 8134 => b:="8134";
                when 8135 => b:="8135";
                when 8136 => b:="8136";
                when 8137 => b:="8137";
                when 8138 => b:="8138";
                when 8139 => b:="8139";
                when 8140 => b:="8140";
                when 8141 => b:="8141";
                when 8142 => b:="8142";
                when 8143 => b:="8143";
                when 8144 => b:="8144";
                when 8145 => b:="8145";
                when 8146 => b:="8146";
                when 8147 => b:="8147";
                when 8148 => b:="8148";
                when 8149 => b:="8149";
                when 8150 => b:="8150";
                when 8151 => b:="8151";
                when 8152 => b:="8152";
                when 8153 => b:="8153";
                when 8154 => b:="8154";
                when 8155 => b:="8155";
                when 8156 => b:="8156";
                when 8157 => b:="8157";
                when 8158 => b:="8158";
                when 8159 => b:="8159";
                when 8160 => b:="8160";
                when 8161 => b:="8161";
                when 8162 => b:="8162";
                when 8163 => b:="8163";
                when 8164 => b:="8164";
                when 8165 => b:="8165";
                when 8166 => b:="8166";
                when 8167 => b:="8167";
                when 8168 => b:="8168";
                when 8169 => b:="8169";
                when 8170 => b:="8170";
                when 8171 => b:="8171";
                when 8172 => b:="8172";
                when 8173 => b:="8173";
                when 8174 => b:="8174";
                when 8175 => b:="8175";
                when 8176 => b:="8176";
                when 8177 => b:="8177";
                when 8178 => b:="8178";
                when 8179 => b:="8179";
                when 8180 => b:="8180";
                when 8181 => b:="8181";
                when 8182 => b:="8182";
                when 8183 => b:="8183";
                when 8184 => b:="8184";
                when 8185 => b:="8185";
                when 8186 => b:="8186";
                when 8187 => b:="8187";
                when 8188 => b:="8188";
                when 8189 => b:="8189";
                when 8190 => b:="8190";
                when 8191 => b:="8191";
                when 8192 => b:="8192";
                when 8193 => b:="8193";
                when 8194 => b:="8194";
                when 8195 => b:="8195";
                when 8196 => b:="8196";
                when 8197 => b:="8197";
                when 8198 => b:="8198";
                when 8199 => b:="8199";
                when 8200 => b:="8200";
                when 8201 => b:="8201";
                when 8202 => b:="8202";
                when 8203 => b:="8203";
                when 8204 => b:="8204";
                when 8205 => b:="8205";
                when 8206 => b:="8206";
                when 8207 => b:="8207";
                when 8208 => b:="8208";
                when 8209 => b:="8209";
                when 8210 => b:="8210";
                when 8211 => b:="8211";
                when 8212 => b:="8212";
                when 8213 => b:="8213";
                when 8214 => b:="8214";
                when 8215 => b:="8215";
                when 8216 => b:="8216";
                when 8217 => b:="8217";
                when 8218 => b:="8218";
                when 8219 => b:="8219";
                when 8220 => b:="8220";
                when 8221 => b:="8221";
                when 8222 => b:="8222";
                when 8223 => b:="8223";
                when 8224 => b:="8224";
                when 8225 => b:="8225";
                when 8226 => b:="8226";
                when 8227 => b:="8227";
                when 8228 => b:="8228";
                when 8229 => b:="8229";
                when 8230 => b:="8230";
                when 8231 => b:="8231";
                when 8232 => b:="8232";
                when 8233 => b:="8233";
                when 8234 => b:="8234";
                when 8235 => b:="8235";
                when 8236 => b:="8236";
                when 8237 => b:="8237";
                when 8238 => b:="8238";
                when 8239 => b:="8239";
                when 8240 => b:="8240";
                when 8241 => b:="8241";
                when 8242 => b:="8242";
                when 8243 => b:="8243";
                when 8244 => b:="8244";
                when 8245 => b:="8245";
                when 8246 => b:="8246";
                when 8247 => b:="8247";
                when 8248 => b:="8248";
                when 8249 => b:="8249";
                when 8250 => b:="8250";
                when 8251 => b:="8251";
                when 8252 => b:="8252";
                when 8253 => b:="8253";
                when 8254 => b:="8254";
                when 8255 => b:="8255";
                when 8256 => b:="8256";
                when 8257 => b:="8257";
                when 8258 => b:="8258";
                when 8259 => b:="8259";
                when 8260 => b:="8260";
                when 8261 => b:="8261";
                when 8262 => b:="8262";
                when 8263 => b:="8263";
                when 8264 => b:="8264";
                when 8265 => b:="8265";
                when 8266 => b:="8266";
                when 8267 => b:="8267";
                when 8268 => b:="8268";
                when 8269 => b:="8269";
                when 8270 => b:="8270";
                when 8271 => b:="8271";
                when 8272 => b:="8272";
                when 8273 => b:="8273";
                when 8274 => b:="8274";
                when 8275 => b:="8275";
                when 8276 => b:="8276";
                when 8277 => b:="8277";
                when 8278 => b:="8278";
                when 8279 => b:="8279";
                when 8280 => b:="8280";
                when 8281 => b:="8281";
                when 8282 => b:="8282";
                when 8283 => b:="8283";
                when 8284 => b:="8284";
                when 8285 => b:="8285";
                when 8286 => b:="8286";
                when 8287 => b:="8287";
                when 8288 => b:="8288";
                when 8289 => b:="8289";
                when 8290 => b:="8290";
                when 8291 => b:="8291";
                when 8292 => b:="8292";
                when 8293 => b:="8293";
                when 8294 => b:="8294";
                when 8295 => b:="8295";
                when 8296 => b:="8296";
                when 8297 => b:="8297";
                when 8298 => b:="8298";
                when 8299 => b:="8299";
                when 8300 => b:="8300";
                when 8301 => b:="8301";
                when 8302 => b:="8302";
                when 8303 => b:="8303";
                when 8304 => b:="8304";
                when 8305 => b:="8305";
                when 8306 => b:="8306";
                when 8307 => b:="8307";
                when 8308 => b:="8308";
                when 8309 => b:="8309";
                when 8310 => b:="8310";
                when 8311 => b:="8311";
                when 8312 => b:="8312";
                when 8313 => b:="8313";
                when 8314 => b:="8314";
                when 8315 => b:="8315";
                when 8316 => b:="8316";
                when 8317 => b:="8317";
                when 8318 => b:="8318";
                when 8319 => b:="8319";
                when 8320 => b:="8320";
                when 8321 => b:="8321";
                when 8322 => b:="8322";
                when 8323 => b:="8323";
                when 8324 => b:="8324";
                when 8325 => b:="8325";
                when 8326 => b:="8326";
                when 8327 => b:="8327";
                when 8328 => b:="8328";
                when 8329 => b:="8329";
                when 8330 => b:="8330";
                when 8331 => b:="8331";
                when 8332 => b:="8332";
                when 8333 => b:="8333";
                when 8334 => b:="8334";
                when 8335 => b:="8335";
                when 8336 => b:="8336";
                when 8337 => b:="8337";
                when 8338 => b:="8338";
                when 8339 => b:="8339";
                when 8340 => b:="8340";
                when 8341 => b:="8341";
                when 8342 => b:="8342";
                when 8343 => b:="8343";
                when 8344 => b:="8344";
                when 8345 => b:="8345";
                when 8346 => b:="8346";
                when 8347 => b:="8347";
                when 8348 => b:="8348";
                when 8349 => b:="8349";
                when 8350 => b:="8350";
                when 8351 => b:="8351";
                when 8352 => b:="8352";
                when 8353 => b:="8353";
                when 8354 => b:="8354";
                when 8355 => b:="8355";
                when 8356 => b:="8356";
                when 8357 => b:="8357";
                when 8358 => b:="8358";
                when 8359 => b:="8359";
                when 8360 => b:="8360";
                when 8361 => b:="8361";
                when 8362 => b:="8362";
                when 8363 => b:="8363";
                when 8364 => b:="8364";
                when 8365 => b:="8365";
                when 8366 => b:="8366";
                when 8367 => b:="8367";
                when 8368 => b:="8368";
                when 8369 => b:="8369";
                when 8370 => b:="8370";
                when 8371 => b:="8371";
                when 8372 => b:="8372";
                when 8373 => b:="8373";
                when 8374 => b:="8374";
                when 8375 => b:="8375";
                when 8376 => b:="8376";
                when 8377 => b:="8377";
                when 8378 => b:="8378";
                when 8379 => b:="8379";
                when 8380 => b:="8380";
                when 8381 => b:="8381";
                when 8382 => b:="8382";
                when 8383 => b:="8383";
                when 8384 => b:="8384";
                when 8385 => b:="8385";
                when 8386 => b:="8386";
                when 8387 => b:="8387";
                when 8388 => b:="8388";
                when 8389 => b:="8389";
                when 8390 => b:="8390";
                when 8391 => b:="8391";
                when 8392 => b:="8392";
                when 8393 => b:="8393";
                when 8394 => b:="8394";
                when 8395 => b:="8395";
                when 8396 => b:="8396";
                when 8397 => b:="8397";
                when 8398 => b:="8398";
                when 8399 => b:="8399";
                when 8400 => b:="8400";
                when 8401 => b:="8401";
                when 8402 => b:="8402";
                when 8403 => b:="8403";
                when 8404 => b:="8404";
                when 8405 => b:="8405";
                when 8406 => b:="8406";
                when 8407 => b:="8407";
                when 8408 => b:="8408";
                when 8409 => b:="8409";
                when 8410 => b:="8410";
                when 8411 => b:="8411";
                when 8412 => b:="8412";
                when 8413 => b:="8413";
                when 8414 => b:="8414";
                when 8415 => b:="8415";
                when 8416 => b:="8416";
                when 8417 => b:="8417";
                when 8418 => b:="8418";
                when 8419 => b:="8419";
                when 8420 => b:="8420";
                when 8421 => b:="8421";
                when 8422 => b:="8422";
                when 8423 => b:="8423";
                when 8424 => b:="8424";
                when 8425 => b:="8425";
                when 8426 => b:="8426";
                when 8427 => b:="8427";
                when 8428 => b:="8428";
                when 8429 => b:="8429";
                when 8430 => b:="8430";
                when 8431 => b:="8431";
                when 8432 => b:="8432";
                when 8433 => b:="8433";
                when 8434 => b:="8434";
                when 8435 => b:="8435";
                when 8436 => b:="8436";
                when 8437 => b:="8437";
                when 8438 => b:="8438";
                when 8439 => b:="8439";
                when 8440 => b:="8440";
                when 8441 => b:="8441";
                when 8442 => b:="8442";
                when 8443 => b:="8443";
                when 8444 => b:="8444";
                when 8445 => b:="8445";
                when 8446 => b:="8446";
                when 8447 => b:="8447";
                when 8448 => b:="8448";
                when 8449 => b:="8449";
                when 8450 => b:="8450";
                when 8451 => b:="8451";
                when 8452 => b:="8452";
                when 8453 => b:="8453";
                when 8454 => b:="8454";
                when 8455 => b:="8455";
                when 8456 => b:="8456";
                when 8457 => b:="8457";
                when 8458 => b:="8458";
                when 8459 => b:="8459";
                when 8460 => b:="8460";
                when 8461 => b:="8461";
                when 8462 => b:="8462";
                when 8463 => b:="8463";
                when 8464 => b:="8464";
                when 8465 => b:="8465";
                when 8466 => b:="8466";
                when 8467 => b:="8467";
                when 8468 => b:="8468";
                when 8469 => b:="8469";
                when 8470 => b:="8470";
                when 8471 => b:="8471";
                when 8472 => b:="8472";
                when 8473 => b:="8473";
                when 8474 => b:="8474";
                when 8475 => b:="8475";
                when 8476 => b:="8476";
                when 8477 => b:="8477";
                when 8478 => b:="8478";
                when 8479 => b:="8479";
                when 8480 => b:="8480";
                when 8481 => b:="8481";
                when 8482 => b:="8482";
                when 8483 => b:="8483";
                when 8484 => b:="8484";
                when 8485 => b:="8485";
                when 8486 => b:="8486";
                when 8487 => b:="8487";
                when 8488 => b:="8488";
                when 8489 => b:="8489";
                when 8490 => b:="8490";
                when 8491 => b:="8491";
                when 8492 => b:="8492";
                when 8493 => b:="8493";
                when 8494 => b:="8494";
                when 8495 => b:="8495";
                when 8496 => b:="8496";
                when 8497 => b:="8497";
                when 8498 => b:="8498";
                when 8499 => b:="8499";
                when 8500 => b:="8500";
                when 8501 => b:="8501";
                when 8502 => b:="8502";
                when 8503 => b:="8503";
                when 8504 => b:="8504";
                when 8505 => b:="8505";
                when 8506 => b:="8506";
                when 8507 => b:="8507";
                when 8508 => b:="8508";
                when 8509 => b:="8509";
                when 8510 => b:="8510";
                when 8511 => b:="8511";
                when 8512 => b:="8512";
                when 8513 => b:="8513";
                when 8514 => b:="8514";
                when 8515 => b:="8515";
                when 8516 => b:="8516";
                when 8517 => b:="8517";
                when 8518 => b:="8518";
                when 8519 => b:="8519";
                when 8520 => b:="8520";
                when 8521 => b:="8521";
                when 8522 => b:="8522";
                when 8523 => b:="8523";
                when 8524 => b:="8524";
                when 8525 => b:="8525";
                when 8526 => b:="8526";
                when 8527 => b:="8527";
                when 8528 => b:="8528";
                when 8529 => b:="8529";
                when 8530 => b:="8530";
                when 8531 => b:="8531";
                when 8532 => b:="8532";
                when 8533 => b:="8533";
                when 8534 => b:="8534";
                when 8535 => b:="8535";
                when 8536 => b:="8536";
                when 8537 => b:="8537";
                when 8538 => b:="8538";
                when 8539 => b:="8539";
                when 8540 => b:="8540";
                when 8541 => b:="8541";
                when 8542 => b:="8542";
                when 8543 => b:="8543";
                when 8544 => b:="8544";
                when 8545 => b:="8545";
                when 8546 => b:="8546";
                when 8547 => b:="8547";
                when 8548 => b:="8548";
                when 8549 => b:="8549";
                when 8550 => b:="8550";
                when 8551 => b:="8551";
                when 8552 => b:="8552";
                when 8553 => b:="8553";
                when 8554 => b:="8554";
                when 8555 => b:="8555";
                when 8556 => b:="8556";
                when 8557 => b:="8557";
                when 8558 => b:="8558";
                when 8559 => b:="8559";
                when 8560 => b:="8560";
                when 8561 => b:="8561";
                when 8562 => b:="8562";
                when 8563 => b:="8563";
                when 8564 => b:="8564";
                when 8565 => b:="8565";
                when 8566 => b:="8566";
                when 8567 => b:="8567";
                when 8568 => b:="8568";
                when 8569 => b:="8569";
                when 8570 => b:="8570";
                when 8571 => b:="8571";
                when 8572 => b:="8572";
                when 8573 => b:="8573";
                when 8574 => b:="8574";
                when 8575 => b:="8575";
                when 8576 => b:="8576";
                when 8577 => b:="8577";
                when 8578 => b:="8578";
                when 8579 => b:="8579";
                when 8580 => b:="8580";
                when 8581 => b:="8581";
                when 8582 => b:="8582";
                when 8583 => b:="8583";
                when 8584 => b:="8584";
                when 8585 => b:="8585";
                when 8586 => b:="8586";
                when 8587 => b:="8587";
                when 8588 => b:="8588";
                when 8589 => b:="8589";
                when 8590 => b:="8590";
                when 8591 => b:="8591";
                when 8592 => b:="8592";
                when 8593 => b:="8593";
                when 8594 => b:="8594";
                when 8595 => b:="8595";
                when 8596 => b:="8596";
                when 8597 => b:="8597";
                when 8598 => b:="8598";
                when 8599 => b:="8599";
                when 8600 => b:="8600";
                when 8601 => b:="8601";
                when 8602 => b:="8602";
                when 8603 => b:="8603";
                when 8604 => b:="8604";
                when 8605 => b:="8605";
                when 8606 => b:="8606";
                when 8607 => b:="8607";
                when 8608 => b:="8608";
                when 8609 => b:="8609";
                when 8610 => b:="8610";
                when 8611 => b:="8611";
                when 8612 => b:="8612";
                when 8613 => b:="8613";
                when 8614 => b:="8614";
                when 8615 => b:="8615";
                when 8616 => b:="8616";
                when 8617 => b:="8617";
                when 8618 => b:="8618";
                when 8619 => b:="8619";
                when 8620 => b:="8620";
                when 8621 => b:="8621";
                when 8622 => b:="8622";
                when 8623 => b:="8623";
                when 8624 => b:="8624";
                when 8625 => b:="8625";
                when 8626 => b:="8626";
                when 8627 => b:="8627";
                when 8628 => b:="8628";
                when 8629 => b:="8629";
                when 8630 => b:="8630";
                when 8631 => b:="8631";
                when 8632 => b:="8632";
                when 8633 => b:="8633";
                when 8634 => b:="8634";
                when 8635 => b:="8635";
                when 8636 => b:="8636";
                when 8637 => b:="8637";
                when 8638 => b:="8638";
                when 8639 => b:="8639";
                when 8640 => b:="8640";
                when 8641 => b:="8641";
                when 8642 => b:="8642";
                when 8643 => b:="8643";
                when 8644 => b:="8644";
                when 8645 => b:="8645";
                when 8646 => b:="8646";
                when 8647 => b:="8647";
                when 8648 => b:="8648";
                when 8649 => b:="8649";
                when 8650 => b:="8650";
                when 8651 => b:="8651";
                when 8652 => b:="8652";
                when 8653 => b:="8653";
                when 8654 => b:="8654";
                when 8655 => b:="8655";
                when 8656 => b:="8656";
                when 8657 => b:="8657";
                when 8658 => b:="8658";
                when 8659 => b:="8659";
                when 8660 => b:="8660";
                when 8661 => b:="8661";
                when 8662 => b:="8662";
                when 8663 => b:="8663";
                when 8664 => b:="8664";
                when 8665 => b:="8665";
                when 8666 => b:="8666";
                when 8667 => b:="8667";
                when 8668 => b:="8668";
                when 8669 => b:="8669";
                when 8670 => b:="8670";
                when 8671 => b:="8671";
                when 8672 => b:="8672";
                when 8673 => b:="8673";
                when 8674 => b:="8674";
                when 8675 => b:="8675";
                when 8676 => b:="8676";
                when 8677 => b:="8677";
                when 8678 => b:="8678";
                when 8679 => b:="8679";
                when 8680 => b:="8680";
                when 8681 => b:="8681";
                when 8682 => b:="8682";
                when 8683 => b:="8683";
                when 8684 => b:="8684";
                when 8685 => b:="8685";
                when 8686 => b:="8686";
                when 8687 => b:="8687";
                when 8688 => b:="8688";
                when 8689 => b:="8689";
                when 8690 => b:="8690";
                when 8691 => b:="8691";
                when 8692 => b:="8692";
                when 8693 => b:="8693";
                when 8694 => b:="8694";
                when 8695 => b:="8695";
                when 8696 => b:="8696";
                when 8697 => b:="8697";
                when 8698 => b:="8698";
                when 8699 => b:="8699";
                when 8700 => b:="8700";
                when 8701 => b:="8701";
                when 8702 => b:="8702";
                when 8703 => b:="8703";
                when 8704 => b:="8704";
                when 8705 => b:="8705";
                when 8706 => b:="8706";
                when 8707 => b:="8707";
                when 8708 => b:="8708";
                when 8709 => b:="8709";
                when 8710 => b:="8710";
                when 8711 => b:="8711";
                when 8712 => b:="8712";
                when 8713 => b:="8713";
                when 8714 => b:="8714";
                when 8715 => b:="8715";
                when 8716 => b:="8716";
                when 8717 => b:="8717";
                when 8718 => b:="8718";
                when 8719 => b:="8719";
                when 8720 => b:="8720";
                when 8721 => b:="8721";
                when 8722 => b:="8722";
                when 8723 => b:="8723";
                when 8724 => b:="8724";
                when 8725 => b:="8725";
                when 8726 => b:="8726";
                when 8727 => b:="8727";
                when 8728 => b:="8728";
                when 8729 => b:="8729";
                when 8730 => b:="8730";
                when 8731 => b:="8731";
                when 8732 => b:="8732";
                when 8733 => b:="8733";
                when 8734 => b:="8734";
                when 8735 => b:="8735";
                when 8736 => b:="8736";
                when 8737 => b:="8737";
                when 8738 => b:="8738";
                when 8739 => b:="8739";
                when 8740 => b:="8740";
                when 8741 => b:="8741";
                when 8742 => b:="8742";
                when 8743 => b:="8743";
                when 8744 => b:="8744";
                when 8745 => b:="8745";
                when 8746 => b:="8746";
                when 8747 => b:="8747";
                when 8748 => b:="8748";
                when 8749 => b:="8749";
                when 8750 => b:="8750";
                when 8751 => b:="8751";
                when 8752 => b:="8752";
                when 8753 => b:="8753";
                when 8754 => b:="8754";
                when 8755 => b:="8755";
                when 8756 => b:="8756";
                when 8757 => b:="8757";
                when 8758 => b:="8758";
                when 8759 => b:="8759";
                when 8760 => b:="8760";
                when 8761 => b:="8761";
                when 8762 => b:="8762";
                when 8763 => b:="8763";
                when 8764 => b:="8764";
                when 8765 => b:="8765";
                when 8766 => b:="8766";
                when 8767 => b:="8767";
                when 8768 => b:="8768";
                when 8769 => b:="8769";
                when 8770 => b:="8770";
                when 8771 => b:="8771";
                when 8772 => b:="8772";
                when 8773 => b:="8773";
                when 8774 => b:="8774";
                when 8775 => b:="8775";
                when 8776 => b:="8776";
                when 8777 => b:="8777";
                when 8778 => b:="8778";
                when 8779 => b:="8779";
                when 8780 => b:="8780";
                when 8781 => b:="8781";
                when 8782 => b:="8782";
                when 8783 => b:="8783";
                when 8784 => b:="8784";
                when 8785 => b:="8785";
                when 8786 => b:="8786";
                when 8787 => b:="8787";
                when 8788 => b:="8788";
                when 8789 => b:="8789";
                when 8790 => b:="8790";
                when 8791 => b:="8791";
                when 8792 => b:="8792";
                when 8793 => b:="8793";
                when 8794 => b:="8794";
                when 8795 => b:="8795";
                when 8796 => b:="8796";
                when 8797 => b:="8797";
                when 8798 => b:="8798";
                when 8799 => b:="8799";
                when 8800 => b:="8800";
                when 8801 => b:="8801";
                when 8802 => b:="8802";
                when 8803 => b:="8803";
                when 8804 => b:="8804";
                when 8805 => b:="8805";
                when 8806 => b:="8806";
                when 8807 => b:="8807";
                when 8808 => b:="8808";
                when 8809 => b:="8809";
                when 8810 => b:="8810";
                when 8811 => b:="8811";
                when 8812 => b:="8812";
                when 8813 => b:="8813";
                when 8814 => b:="8814";
                when 8815 => b:="8815";
                when 8816 => b:="8816";
                when 8817 => b:="8817";
                when 8818 => b:="8818";
                when 8819 => b:="8819";
                when 8820 => b:="8820";
                when 8821 => b:="8821";
                when 8822 => b:="8822";
                when 8823 => b:="8823";
                when 8824 => b:="8824";
                when 8825 => b:="8825";
                when 8826 => b:="8826";
                when 8827 => b:="8827";
                when 8828 => b:="8828";
                when 8829 => b:="8829";
                when 8830 => b:="8830";
                when 8831 => b:="8831";
                when 8832 => b:="8832";
                when 8833 => b:="8833";
                when 8834 => b:="8834";
                when 8835 => b:="8835";
                when 8836 => b:="8836";
                when 8837 => b:="8837";
                when 8838 => b:="8838";
                when 8839 => b:="8839";
                when 8840 => b:="8840";
                when 8841 => b:="8841";
                when 8842 => b:="8842";
                when 8843 => b:="8843";
                when 8844 => b:="8844";
                when 8845 => b:="8845";
                when 8846 => b:="8846";
                when 8847 => b:="8847";
                when 8848 => b:="8848";
                when 8849 => b:="8849";
                when 8850 => b:="8850";
                when 8851 => b:="8851";
                when 8852 => b:="8852";
                when 8853 => b:="8853";
                when 8854 => b:="8854";
                when 8855 => b:="8855";
                when 8856 => b:="8856";
                when 8857 => b:="8857";
                when 8858 => b:="8858";
                when 8859 => b:="8859";
                when 8860 => b:="8860";
                when 8861 => b:="8861";
                when 8862 => b:="8862";
                when 8863 => b:="8863";
                when 8864 => b:="8864";
                when 8865 => b:="8865";
                when 8866 => b:="8866";
                when 8867 => b:="8867";
                when 8868 => b:="8868";
                when 8869 => b:="8869";
                when 8870 => b:="8870";
                when 8871 => b:="8871";
                when 8872 => b:="8872";
                when 8873 => b:="8873";
                when 8874 => b:="8874";
                when 8875 => b:="8875";
                when 8876 => b:="8876";
                when 8877 => b:="8877";
                when 8878 => b:="8878";
                when 8879 => b:="8879";
                when 8880 => b:="8880";
                when 8881 => b:="8881";
                when 8882 => b:="8882";
                when 8883 => b:="8883";
                when 8884 => b:="8884";
                when 8885 => b:="8885";
                when 8886 => b:="8886";
                when 8887 => b:="8887";
                when 8888 => b:="8888";
                when 8889 => b:="8889";
                when 8890 => b:="8890";
                when 8891 => b:="8891";
                when 8892 => b:="8892";
                when 8893 => b:="8893";
                when 8894 => b:="8894";
                when 8895 => b:="8895";
                when 8896 => b:="8896";
                when 8897 => b:="8897";
                when 8898 => b:="8898";
                when 8899 => b:="8899";
                when 8900 => b:="8900";
                when 8901 => b:="8901";
                when 8902 => b:="8902";
                when 8903 => b:="8903";
                when 8904 => b:="8904";
                when 8905 => b:="8905";
                when 8906 => b:="8906";
                when 8907 => b:="8907";
                when 8908 => b:="8908";
                when 8909 => b:="8909";
                when 8910 => b:="8910";
                when 8911 => b:="8911";
                when 8912 => b:="8912";
                when 8913 => b:="8913";
                when 8914 => b:="8914";
                when 8915 => b:="8915";
                when 8916 => b:="8916";
                when 8917 => b:="8917";
                when 8918 => b:="8918";
                when 8919 => b:="8919";
                when 8920 => b:="8920";
                when 8921 => b:="8921";
                when 8922 => b:="8922";
                when 8923 => b:="8923";
                when 8924 => b:="8924";
                when 8925 => b:="8925";
                when 8926 => b:="8926";
                when 8927 => b:="8927";
                when 8928 => b:="8928";
                when 8929 => b:="8929";
                when 8930 => b:="8930";
                when 8931 => b:="8931";
                when 8932 => b:="8932";
                when 8933 => b:="8933";
                when 8934 => b:="8934";
                when 8935 => b:="8935";
                when 8936 => b:="8936";
                when 8937 => b:="8937";
                when 8938 => b:="8938";
                when 8939 => b:="8939";
                when 8940 => b:="8940";
                when 8941 => b:="8941";
                when 8942 => b:="8942";
                when 8943 => b:="8943";
                when 8944 => b:="8944";
                when 8945 => b:="8945";
                when 8946 => b:="8946";
                when 8947 => b:="8947";
                when 8948 => b:="8948";
                when 8949 => b:="8949";
                when 8950 => b:="8950";
                when 8951 => b:="8951";
                when 8952 => b:="8952";
                when 8953 => b:="8953";
                when 8954 => b:="8954";
                when 8955 => b:="8955";
                when 8956 => b:="8956";
                when 8957 => b:="8957";
                when 8958 => b:="8958";
                when 8959 => b:="8959";
                when 8960 => b:="8960";
                when 8961 => b:="8961";
                when 8962 => b:="8962";
                when 8963 => b:="8963";
                when 8964 => b:="8964";
                when 8965 => b:="8965";
                when 8966 => b:="8966";
                when 8967 => b:="8967";
                when 8968 => b:="8968";
                when 8969 => b:="8969";
                when 8970 => b:="8970";
                when 8971 => b:="8971";
                when 8972 => b:="8972";
                when 8973 => b:="8973";
                when 8974 => b:="8974";
                when 8975 => b:="8975";
                when 8976 => b:="8976";
                when 8977 => b:="8977";
                when 8978 => b:="8978";
                when 8979 => b:="8979";
                when 8980 => b:="8980";
                when 8981 => b:="8981";
                when 8982 => b:="8982";
                when 8983 => b:="8983";
                when 8984 => b:="8984";
                when 8985 => b:="8985";
                when 8986 => b:="8986";
                when 8987 => b:="8987";
                when 8988 => b:="8988";
                when 8989 => b:="8989";
                when 8990 => b:="8990";
                when 8991 => b:="8991";
                when 8992 => b:="8992";
                when 8993 => b:="8993";
                when 8994 => b:="8994";
                when 8995 => b:="8995";
                when 8996 => b:="8996";
                when 8997 => b:="8997";
                when 8998 => b:="8998";
                when 8999 => b:="8999";
                when 9000 => b:="9000";
                when 9001 => b:="9001";
                when 9002 => b:="9002";
                when 9003 => b:="9003";
                when 9004 => b:="9004";
                when 9005 => b:="9005";
                when 9006 => b:="9006";
                when 9007 => b:="9007";
                when 9008 => b:="9008";
                when 9009 => b:="9009";
                when 9010 => b:="9010";
                when 9011 => b:="9011";
                when 9012 => b:="9012";
                when 9013 => b:="9013";
                when 9014 => b:="9014";
                when 9015 => b:="9015";
                when 9016 => b:="9016";
                when 9017 => b:="9017";
                when 9018 => b:="9018";
                when 9019 => b:="9019";
                when 9020 => b:="9020";
                when 9021 => b:="9021";
                when 9022 => b:="9022";
                when 9023 => b:="9023";
                when 9024 => b:="9024";
                when 9025 => b:="9025";
                when 9026 => b:="9026";
                when 9027 => b:="9027";
                when 9028 => b:="9028";
                when 9029 => b:="9029";
                when 9030 => b:="9030";
                when 9031 => b:="9031";
                when 9032 => b:="9032";
                when 9033 => b:="9033";
                when 9034 => b:="9034";
                when 9035 => b:="9035";
                when 9036 => b:="9036";
                when 9037 => b:="9037";
                when 9038 => b:="9038";
                when 9039 => b:="9039";
                when 9040 => b:="9040";
                when 9041 => b:="9041";
                when 9042 => b:="9042";
                when 9043 => b:="9043";
                when 9044 => b:="9044";
                when 9045 => b:="9045";
                when 9046 => b:="9046";
                when 9047 => b:="9047";
                when 9048 => b:="9048";
                when 9049 => b:="9049";
                when 9050 => b:="9050";
                when 9051 => b:="9051";
                when 9052 => b:="9052";
                when 9053 => b:="9053";
                when 9054 => b:="9054";
                when 9055 => b:="9055";
                when 9056 => b:="9056";
                when 9057 => b:="9057";
                when 9058 => b:="9058";
                when 9059 => b:="9059";
                when 9060 => b:="9060";
                when 9061 => b:="9061";
                when 9062 => b:="9062";
                when 9063 => b:="9063";
                when 9064 => b:="9064";
                when 9065 => b:="9065";
                when 9066 => b:="9066";
                when 9067 => b:="9067";
                when 9068 => b:="9068";
                when 9069 => b:="9069";
                when 9070 => b:="9070";
                when 9071 => b:="9071";
                when 9072 => b:="9072";
                when 9073 => b:="9073";
                when 9074 => b:="9074";
                when 9075 => b:="9075";
                when 9076 => b:="9076";
                when 9077 => b:="9077";
                when 9078 => b:="9078";
                when 9079 => b:="9079";
                when 9080 => b:="9080";
                when 9081 => b:="9081";
                when 9082 => b:="9082";
                when 9083 => b:="9083";
                when 9084 => b:="9084";
                when 9085 => b:="9085";
                when 9086 => b:="9086";
                when 9087 => b:="9087";
                when 9088 => b:="9088";
                when 9089 => b:="9089";
                when 9090 => b:="9090";
                when 9091 => b:="9091";
                when 9092 => b:="9092";
                when 9093 => b:="9093";
                when 9094 => b:="9094";
                when 9095 => b:="9095";
                when 9096 => b:="9096";
                when 9097 => b:="9097";
                when 9098 => b:="9098";
                when 9099 => b:="9099";
                when 9100 => b:="9100";
                when 9101 => b:="9101";
                when 9102 => b:="9102";
                when 9103 => b:="9103";
                when 9104 => b:="9104";
                when 9105 => b:="9105";
                when 9106 => b:="9106";
                when 9107 => b:="9107";
                when 9108 => b:="9108";
                when 9109 => b:="9109";
                when 9110 => b:="9110";
                when 9111 => b:="9111";
                when 9112 => b:="9112";
                when 9113 => b:="9113";
                when 9114 => b:="9114";
                when 9115 => b:="9115";
                when 9116 => b:="9116";
                when 9117 => b:="9117";
                when 9118 => b:="9118";
                when 9119 => b:="9119";
                when 9120 => b:="9120";
                when 9121 => b:="9121";
                when 9122 => b:="9122";
                when 9123 => b:="9123";
                when 9124 => b:="9124";
                when 9125 => b:="9125";
                when 9126 => b:="9126";
                when 9127 => b:="9127";
                when 9128 => b:="9128";
                when 9129 => b:="9129";
                when 9130 => b:="9130";
                when 9131 => b:="9131";
                when 9132 => b:="9132";
                when 9133 => b:="9133";
                when 9134 => b:="9134";
                when 9135 => b:="9135";
                when 9136 => b:="9136";
                when 9137 => b:="9137";
                when 9138 => b:="9138";
                when 9139 => b:="9139";
                when 9140 => b:="9140";
                when 9141 => b:="9141";
                when 9142 => b:="9142";
                when 9143 => b:="9143";
                when 9144 => b:="9144";
                when 9145 => b:="9145";
                when 9146 => b:="9146";
                when 9147 => b:="9147";
                when 9148 => b:="9148";
                when 9149 => b:="9149";
                when 9150 => b:="9150";
                when 9151 => b:="9151";
                when 9152 => b:="9152";
                when 9153 => b:="9153";
                when 9154 => b:="9154";
                when 9155 => b:="9155";
                when 9156 => b:="9156";
                when 9157 => b:="9157";
                when 9158 => b:="9158";
                when 9159 => b:="9159";
                when 9160 => b:="9160";
                when 9161 => b:="9161";
                when 9162 => b:="9162";
                when 9163 => b:="9163";
                when 9164 => b:="9164";
                when 9165 => b:="9165";
                when 9166 => b:="9166";
                when 9167 => b:="9167";
                when 9168 => b:="9168";
                when 9169 => b:="9169";
                when 9170 => b:="9170";
                when 9171 => b:="9171";
                when 9172 => b:="9172";
                when 9173 => b:="9173";
                when 9174 => b:="9174";
                when 9175 => b:="9175";
                when 9176 => b:="9176";
                when 9177 => b:="9177";
                when 9178 => b:="9178";
                when 9179 => b:="9179";
                when 9180 => b:="9180";
                when 9181 => b:="9181";
                when 9182 => b:="9182";
                when 9183 => b:="9183";
                when 9184 => b:="9184";
                when 9185 => b:="9185";
                when 9186 => b:="9186";
                when 9187 => b:="9187";
                when 9188 => b:="9188";
                when 9189 => b:="9189";
                when 9190 => b:="9190";
                when 9191 => b:="9191";
                when 9192 => b:="9192";
                when 9193 => b:="9193";
                when 9194 => b:="9194";
                when 9195 => b:="9195";
                when 9196 => b:="9196";
                when 9197 => b:="9197";
                when 9198 => b:="9198";
                when 9199 => b:="9199";
                when 9200 => b:="9200";
                when 9201 => b:="9201";
                when 9202 => b:="9202";
                when 9203 => b:="9203";
                when 9204 => b:="9204";
                when 9205 => b:="9205";
                when 9206 => b:="9206";
                when 9207 => b:="9207";
                when 9208 => b:="9208";
                when 9209 => b:="9209";
                when 9210 => b:="9210";
                when 9211 => b:="9211";
                when 9212 => b:="9212";
                when 9213 => b:="9213";
                when 9214 => b:="9214";
                when 9215 => b:="9215";
                when 9216 => b:="9216";
                when 9217 => b:="9217";
                when 9218 => b:="9218";
                when 9219 => b:="9219";
                when 9220 => b:="9220";
                when 9221 => b:="9221";
                when 9222 => b:="9222";
                when 9223 => b:="9223";
                when 9224 => b:="9224";
                when 9225 => b:="9225";
                when 9226 => b:="9226";
                when 9227 => b:="9227";
                when 9228 => b:="9228";
                when 9229 => b:="9229";
                when 9230 => b:="9230";
                when 9231 => b:="9231";
                when 9232 => b:="9232";
                when 9233 => b:="9233";
                when 9234 => b:="9234";
                when 9235 => b:="9235";
                when 9236 => b:="9236";
                when 9237 => b:="9237";
                when 9238 => b:="9238";
                when 9239 => b:="9239";
                when 9240 => b:="9240";
                when 9241 => b:="9241";
                when 9242 => b:="9242";
                when 9243 => b:="9243";
                when 9244 => b:="9244";
                when 9245 => b:="9245";
                when 9246 => b:="9246";
                when 9247 => b:="9247";
                when 9248 => b:="9248";
                when 9249 => b:="9249";
                when 9250 => b:="9250";
                when 9251 => b:="9251";
                when 9252 => b:="9252";
                when 9253 => b:="9253";
                when 9254 => b:="9254";
                when 9255 => b:="9255";
                when 9256 => b:="9256";
                when 9257 => b:="9257";
                when 9258 => b:="9258";
                when 9259 => b:="9259";
                when 9260 => b:="9260";
                when 9261 => b:="9261";
                when 9262 => b:="9262";
                when 9263 => b:="9263";
                when 9264 => b:="9264";
                when 9265 => b:="9265";
                when 9266 => b:="9266";
                when 9267 => b:="9267";
                when 9268 => b:="9268";
                when 9269 => b:="9269";
                when 9270 => b:="9270";
                when 9271 => b:="9271";
                when 9272 => b:="9272";
                when 9273 => b:="9273";
                when 9274 => b:="9274";
                when 9275 => b:="9275";
                when 9276 => b:="9276";
                when 9277 => b:="9277";
                when 9278 => b:="9278";
                when 9279 => b:="9279";
                when 9280 => b:="9280";
                when 9281 => b:="9281";
                when 9282 => b:="9282";
                when 9283 => b:="9283";
                when 9284 => b:="9284";
                when 9285 => b:="9285";
                when 9286 => b:="9286";
                when 9287 => b:="9287";
                when 9288 => b:="9288";
                when 9289 => b:="9289";
                when 9290 => b:="9290";
                when 9291 => b:="9291";
                when 9292 => b:="9292";
                when 9293 => b:="9293";
                when 9294 => b:="9294";
                when 9295 => b:="9295";
                when 9296 => b:="9296";
                when 9297 => b:="9297";
                when 9298 => b:="9298";
                when 9299 => b:="9299";
                when 9300 => b:="9300";
                when 9301 => b:="9301";
                when 9302 => b:="9302";
                when 9303 => b:="9303";
                when 9304 => b:="9304";
                when 9305 => b:="9305";
                when 9306 => b:="9306";
                when 9307 => b:="9307";
                when 9308 => b:="9308";
                when 9309 => b:="9309";
                when 9310 => b:="9310";
                when 9311 => b:="9311";
                when 9312 => b:="9312";
                when 9313 => b:="9313";
                when 9314 => b:="9314";
                when 9315 => b:="9315";
                when 9316 => b:="9316";
                when 9317 => b:="9317";
                when 9318 => b:="9318";
                when 9319 => b:="9319";
                when 9320 => b:="9320";
                when 9321 => b:="9321";
                when 9322 => b:="9322";
                when 9323 => b:="9323";
                when 9324 => b:="9324";
                when 9325 => b:="9325";
                when 9326 => b:="9326";
                when 9327 => b:="9327";
                when 9328 => b:="9328";
                when 9329 => b:="9329";
                when 9330 => b:="9330";
                when 9331 => b:="9331";
                when 9332 => b:="9332";
                when 9333 => b:="9333";
                when 9334 => b:="9334";
                when 9335 => b:="9335";
                when 9336 => b:="9336";
                when 9337 => b:="9337";
                when 9338 => b:="9338";
                when 9339 => b:="9339";
                when 9340 => b:="9340";
                when 9341 => b:="9341";
                when 9342 => b:="9342";
                when 9343 => b:="9343";
                when 9344 => b:="9344";
                when 9345 => b:="9345";
                when 9346 => b:="9346";
                when 9347 => b:="9347";
                when 9348 => b:="9348";
                when 9349 => b:="9349";
                when 9350 => b:="9350";
                when 9351 => b:="9351";
                when 9352 => b:="9352";
                when 9353 => b:="9353";
                when 9354 => b:="9354";
                when 9355 => b:="9355";
                when 9356 => b:="9356";
                when 9357 => b:="9357";
                when 9358 => b:="9358";
                when 9359 => b:="9359";
                when 9360 => b:="9360";
                when 9361 => b:="9361";
                when 9362 => b:="9362";
                when 9363 => b:="9363";
                when 9364 => b:="9364";
                when 9365 => b:="9365";
                when 9366 => b:="9366";
                when 9367 => b:="9367";
                when 9368 => b:="9368";
                when 9369 => b:="9369";
                when 9370 => b:="9370";
                when 9371 => b:="9371";
                when 9372 => b:="9372";
                when 9373 => b:="9373";
                when 9374 => b:="9374";
                when 9375 => b:="9375";
                when 9376 => b:="9376";
                when 9377 => b:="9377";
                when 9378 => b:="9378";
                when 9379 => b:="9379";
                when 9380 => b:="9380";
                when 9381 => b:="9381";
                when 9382 => b:="9382";
                when 9383 => b:="9383";
                when 9384 => b:="9384";
                when 9385 => b:="9385";
                when 9386 => b:="9386";
                when 9387 => b:="9387";
                when 9388 => b:="9388";
                when 9389 => b:="9389";
                when 9390 => b:="9390";
                when 9391 => b:="9391";
                when 9392 => b:="9392";
                when 9393 => b:="9393";
                when 9394 => b:="9394";
                when 9395 => b:="9395";
                when 9396 => b:="9396";
                when 9397 => b:="9397";
                when 9398 => b:="9398";
                when 9399 => b:="9399";
                when 9400 => b:="9400";
                when 9401 => b:="9401";
                when 9402 => b:="9402";
                when 9403 => b:="9403";
                when 9404 => b:="9404";
                when 9405 => b:="9405";
                when 9406 => b:="9406";
                when 9407 => b:="9407";
                when 9408 => b:="9408";
                when 9409 => b:="9409";
                when 9410 => b:="9410";
                when 9411 => b:="9411";
                when 9412 => b:="9412";
                when 9413 => b:="9413";
                when 9414 => b:="9414";
                when 9415 => b:="9415";
                when 9416 => b:="9416";
                when 9417 => b:="9417";
                when 9418 => b:="9418";
                when 9419 => b:="9419";
                when 9420 => b:="9420";
                when 9421 => b:="9421";
                when 9422 => b:="9422";
                when 9423 => b:="9423";
                when 9424 => b:="9424";
                when 9425 => b:="9425";
                when 9426 => b:="9426";
                when 9427 => b:="9427";
                when 9428 => b:="9428";
                when 9429 => b:="9429";
                when 9430 => b:="9430";
                when 9431 => b:="9431";
                when 9432 => b:="9432";
                when 9433 => b:="9433";
                when 9434 => b:="9434";
                when 9435 => b:="9435";
                when 9436 => b:="9436";
                when 9437 => b:="9437";
                when 9438 => b:="9438";
                when 9439 => b:="9439";
                when 9440 => b:="9440";
                when 9441 => b:="9441";
                when 9442 => b:="9442";
                when 9443 => b:="9443";
                when 9444 => b:="9444";
                when 9445 => b:="9445";
                when 9446 => b:="9446";
                when 9447 => b:="9447";
                when 9448 => b:="9448";
                when 9449 => b:="9449";
                when 9450 => b:="9450";
                when 9451 => b:="9451";
                when 9452 => b:="9452";
                when 9453 => b:="9453";
                when 9454 => b:="9454";
                when 9455 => b:="9455";
                when 9456 => b:="9456";
                when 9457 => b:="9457";
                when 9458 => b:="9458";
                when 9459 => b:="9459";
                when 9460 => b:="9460";
                when 9461 => b:="9461";
                when 9462 => b:="9462";
                when 9463 => b:="9463";
                when 9464 => b:="9464";
                when 9465 => b:="9465";
                when 9466 => b:="9466";
                when 9467 => b:="9467";
                when 9468 => b:="9468";
                when 9469 => b:="9469";
                when 9470 => b:="9470";
                when 9471 => b:="9471";
                when 9472 => b:="9472";
                when 9473 => b:="9473";
                when 9474 => b:="9474";
                when 9475 => b:="9475";
                when 9476 => b:="9476";
                when 9477 => b:="9477";
                when 9478 => b:="9478";
                when 9479 => b:="9479";
                when 9480 => b:="9480";
                when 9481 => b:="9481";
                when 9482 => b:="9482";
                when 9483 => b:="9483";
                when 9484 => b:="9484";
                when 9485 => b:="9485";
                when 9486 => b:="9486";
                when 9487 => b:="9487";
                when 9488 => b:="9488";
                when 9489 => b:="9489";
                when 9490 => b:="9490";
                when 9491 => b:="9491";
                when 9492 => b:="9492";
                when 9493 => b:="9493";
                when 9494 => b:="9494";
                when 9495 => b:="9495";
                when 9496 => b:="9496";
                when 9497 => b:="9497";
                when 9498 => b:="9498";
                when 9499 => b:="9499";
                when 9500 => b:="9500";
                when 9501 => b:="9501";
                when 9502 => b:="9502";
                when 9503 => b:="9503";
                when 9504 => b:="9504";
                when 9505 => b:="9505";
                when 9506 => b:="9506";
                when 9507 => b:="9507";
                when 9508 => b:="9508";
                when 9509 => b:="9509";
                when 9510 => b:="9510";
                when 9511 => b:="9511";
                when 9512 => b:="9512";
                when 9513 => b:="9513";
                when 9514 => b:="9514";
                when 9515 => b:="9515";
                when 9516 => b:="9516";
                when 9517 => b:="9517";
                when 9518 => b:="9518";
                when 9519 => b:="9519";
                when 9520 => b:="9520";
                when 9521 => b:="9521";
                when 9522 => b:="9522";
                when 9523 => b:="9523";
                when 9524 => b:="9524";
                when 9525 => b:="9525";
                when 9526 => b:="9526";
                when 9527 => b:="9527";
                when 9528 => b:="9528";
                when 9529 => b:="9529";
                when 9530 => b:="9530";
                when 9531 => b:="9531";
                when 9532 => b:="9532";
                when 9533 => b:="9533";
                when 9534 => b:="9534";
                when 9535 => b:="9535";
                when 9536 => b:="9536";
                when 9537 => b:="9537";
                when 9538 => b:="9538";
                when 9539 => b:="9539";
                when 9540 => b:="9540";
                when 9541 => b:="9541";
                when 9542 => b:="9542";
                when 9543 => b:="9543";
                when 9544 => b:="9544";
                when 9545 => b:="9545";
                when 9546 => b:="9546";
                when 9547 => b:="9547";
                when 9548 => b:="9548";
                when 9549 => b:="9549";
                when 9550 => b:="9550";
                when 9551 => b:="9551";
                when 9552 => b:="9552";
                when 9553 => b:="9553";
                when 9554 => b:="9554";
                when 9555 => b:="9555";
                when 9556 => b:="9556";
                when 9557 => b:="9557";
                when 9558 => b:="9558";
                when 9559 => b:="9559";
                when 9560 => b:="9560";
                when 9561 => b:="9561";
                when 9562 => b:="9562";
                when 9563 => b:="9563";
                when 9564 => b:="9564";
                when 9565 => b:="9565";
                when 9566 => b:="9566";
                when 9567 => b:="9567";
                when 9568 => b:="9568";
                when 9569 => b:="9569";
                when 9570 => b:="9570";
                when 9571 => b:="9571";
                when 9572 => b:="9572";
                when 9573 => b:="9573";
                when 9574 => b:="9574";
                when 9575 => b:="9575";
                when 9576 => b:="9576";
                when 9577 => b:="9577";
                when 9578 => b:="9578";
                when 9579 => b:="9579";
                when 9580 => b:="9580";
                when 9581 => b:="9581";
                when 9582 => b:="9582";
                when 9583 => b:="9583";
                when 9584 => b:="9584";
                when 9585 => b:="9585";
                when 9586 => b:="9586";
                when 9587 => b:="9587";
                when 9588 => b:="9588";
                when 9589 => b:="9589";
                when 9590 => b:="9590";
                when 9591 => b:="9591";
                when 9592 => b:="9592";
                when 9593 => b:="9593";
                when 9594 => b:="9594";
                when 9595 => b:="9595";
                when 9596 => b:="9596";
                when 9597 => b:="9597";
                when 9598 => b:="9598";
                when 9599 => b:="9599";
                when 9600 => b:="9600";
                when 9601 => b:="9601";
                when 9602 => b:="9602";
                when 9603 => b:="9603";
                when 9604 => b:="9604";
                when 9605 => b:="9605";
                when 9606 => b:="9606";
                when 9607 => b:="9607";
                when 9608 => b:="9608";
                when 9609 => b:="9609";
                when 9610 => b:="9610";
                when 9611 => b:="9611";
                when 9612 => b:="9612";
                when 9613 => b:="9613";
                when 9614 => b:="9614";
                when 9615 => b:="9615";
                when 9616 => b:="9616";
                when 9617 => b:="9617";
                when 9618 => b:="9618";
                when 9619 => b:="9619";
                when 9620 => b:="9620";
                when 9621 => b:="9621";
                when 9622 => b:="9622";
                when 9623 => b:="9623";
                when 9624 => b:="9624";
                when 9625 => b:="9625";
                when 9626 => b:="9626";
                when 9627 => b:="9627";
                when 9628 => b:="9628";
                when 9629 => b:="9629";
                when 9630 => b:="9630";
                when 9631 => b:="9631";
                when 9632 => b:="9632";
                when 9633 => b:="9633";
                when 9634 => b:="9634";
                when 9635 => b:="9635";
                when 9636 => b:="9636";
                when 9637 => b:="9637";
                when 9638 => b:="9638";
                when 9639 => b:="9639";
                when 9640 => b:="9640";
                when 9641 => b:="9641";
                when 9642 => b:="9642";
                when 9643 => b:="9643";
                when 9644 => b:="9644";
                when 9645 => b:="9645";
                when 9646 => b:="9646";
                when 9647 => b:="9647";
                when 9648 => b:="9648";
                when 9649 => b:="9649";
                when 9650 => b:="9650";
                when 9651 => b:="9651";
                when 9652 => b:="9652";
                when 9653 => b:="9653";
                when 9654 => b:="9654";
                when 9655 => b:="9655";
                when 9656 => b:="9656";
                when 9657 => b:="9657";
                when 9658 => b:="9658";
                when 9659 => b:="9659";
                when 9660 => b:="9660";
                when 9661 => b:="9661";
                when 9662 => b:="9662";
                when 9663 => b:="9663";
                when 9664 => b:="9664";
                when 9665 => b:="9665";
                when 9666 => b:="9666";
                when 9667 => b:="9667";
                when 9668 => b:="9668";
                when 9669 => b:="9669";
                when 9670 => b:="9670";
                when 9671 => b:="9671";
                when 9672 => b:="9672";
                when 9673 => b:="9673";
                when 9674 => b:="9674";
                when 9675 => b:="9675";
                when 9676 => b:="9676";
                when 9677 => b:="9677";
                when 9678 => b:="9678";
                when 9679 => b:="9679";
                when 9680 => b:="9680";
                when 9681 => b:="9681";
                when 9682 => b:="9682";
                when 9683 => b:="9683";
                when 9684 => b:="9684";
                when 9685 => b:="9685";
                when 9686 => b:="9686";
                when 9687 => b:="9687";
                when 9688 => b:="9688";
                when 9689 => b:="9689";
                when 9690 => b:="9690";
                when 9691 => b:="9691";
                when 9692 => b:="9692";
                when 9693 => b:="9693";
                when 9694 => b:="9694";
                when 9695 => b:="9695";
                when 9696 => b:="9696";
                when 9697 => b:="9697";
                when 9698 => b:="9698";
                when 9699 => b:="9699";
                when 9700 => b:="9700";
                when 9701 => b:="9701";
                when 9702 => b:="9702";
                when 9703 => b:="9703";
                when 9704 => b:="9704";
                when 9705 => b:="9705";
                when 9706 => b:="9706";
                when 9707 => b:="9707";
                when 9708 => b:="9708";
                when 9709 => b:="9709";
                when 9710 => b:="9710";
                when 9711 => b:="9711";
                when 9712 => b:="9712";
                when 9713 => b:="9713";
                when 9714 => b:="9714";
                when 9715 => b:="9715";
                when 9716 => b:="9716";
                when 9717 => b:="9717";
                when 9718 => b:="9718";
                when 9719 => b:="9719";
                when 9720 => b:="9720";
                when 9721 => b:="9721";
                when 9722 => b:="9722";
                when 9723 => b:="9723";
                when 9724 => b:="9724";
                when 9725 => b:="9725";
                when 9726 => b:="9726";
                when 9727 => b:="9727";
                when 9728 => b:="9728";
                when 9729 => b:="9729";
                when 9730 => b:="9730";
                when 9731 => b:="9731";
                when 9732 => b:="9732";
                when 9733 => b:="9733";
                when 9734 => b:="9734";
                when 9735 => b:="9735";
                when 9736 => b:="9736";
                when 9737 => b:="9737";
                when 9738 => b:="9738";
                when 9739 => b:="9739";
                when 9740 => b:="9740";
                when 9741 => b:="9741";
                when 9742 => b:="9742";
                when 9743 => b:="9743";
                when 9744 => b:="9744";
                when 9745 => b:="9745";
                when 9746 => b:="9746";
                when 9747 => b:="9747";
                when 9748 => b:="9748";
                when 9749 => b:="9749";
                when 9750 => b:="9750";
                when 9751 => b:="9751";
                when 9752 => b:="9752";
                when 9753 => b:="9753";
                when 9754 => b:="9754";
                when 9755 => b:="9755";
                when 9756 => b:="9756";
                when 9757 => b:="9757";
                when 9758 => b:="9758";
                when 9759 => b:="9759";
                when 9760 => b:="9760";
                when 9761 => b:="9761";
                when 9762 => b:="9762";
                when 9763 => b:="9763";
                when 9764 => b:="9764";
                when 9765 => b:="9765";
                when 9766 => b:="9766";
                when 9767 => b:="9767";
                when 9768 => b:="9768";
                when 9769 => b:="9769";
                when 9770 => b:="9770";
                when 9771 => b:="9771";
                when 9772 => b:="9772";
                when 9773 => b:="9773";
                when 9774 => b:="9774";
                when 9775 => b:="9775";
                when 9776 => b:="9776";
                when 9777 => b:="9777";
                when 9778 => b:="9778";
                when 9779 => b:="9779";
                when 9780 => b:="9780";
                when 9781 => b:="9781";
                when 9782 => b:="9782";
                when 9783 => b:="9783";
                when 9784 => b:="9784";
                when 9785 => b:="9785";
                when 9786 => b:="9786";
                when 9787 => b:="9787";
                when 9788 => b:="9788";
                when 9789 => b:="9789";
                when 9790 => b:="9790";
                when 9791 => b:="9791";
                when 9792 => b:="9792";
                when 9793 => b:="9793";
                when 9794 => b:="9794";
                when 9795 => b:="9795";
                when 9796 => b:="9796";
                when 9797 => b:="9797";
                when 9798 => b:="9798";
                when 9799 => b:="9799";
                when 9800 => b:="9800";
                when 9801 => b:="9801";
                when 9802 => b:="9802";
                when 9803 => b:="9803";
                when 9804 => b:="9804";
                when 9805 => b:="9805";
                when 9806 => b:="9806";
                when 9807 => b:="9807";
                when 9808 => b:="9808";
                when 9809 => b:="9809";
                when 9810 => b:="9810";
                when 9811 => b:="9811";
                when 9812 => b:="9812";
                when 9813 => b:="9813";
                when 9814 => b:="9814";
                when 9815 => b:="9815";
                when 9816 => b:="9816";
                when 9817 => b:="9817";
                when 9818 => b:="9818";
                when 9819 => b:="9819";
                when 9820 => b:="9820";
                when 9821 => b:="9821";
                when 9822 => b:="9822";
                when 9823 => b:="9823";
                when 9824 => b:="9824";
                when 9825 => b:="9825";
                when 9826 => b:="9826";
                when 9827 => b:="9827";
                when 9828 => b:="9828";
                when 9829 => b:="9829";
                when 9830 => b:="9830";
                when 9831 => b:="9831";
                when 9832 => b:="9832";
                when 9833 => b:="9833";
                when 9834 => b:="9834";
                when 9835 => b:="9835";
                when 9836 => b:="9836";
                when 9837 => b:="9837";
                when 9838 => b:="9838";
                when 9839 => b:="9839";
                when 9840 => b:="9840";
                when 9841 => b:="9841";
                when 9842 => b:="9842";
                when 9843 => b:="9843";
                when 9844 => b:="9844";
                when 9845 => b:="9845";
                when 9846 => b:="9846";
                when 9847 => b:="9847";
                when 9848 => b:="9848";
                when 9849 => b:="9849";
                when 9850 => b:="9850";
                when 9851 => b:="9851";
                when 9852 => b:="9852";
                when 9853 => b:="9853";
                when 9854 => b:="9854";
                when 9855 => b:="9855";
                when 9856 => b:="9856";
                when 9857 => b:="9857";
                when 9858 => b:="9858";
                when 9859 => b:="9859";
                when 9860 => b:="9860";
                when 9861 => b:="9861";
                when 9862 => b:="9862";
                when 9863 => b:="9863";
                when 9864 => b:="9864";
                when 9865 => b:="9865";
                when 9866 => b:="9866";
                when 9867 => b:="9867";
                when 9868 => b:="9868";
                when 9869 => b:="9869";
                when 9870 => b:="9870";
                when 9871 => b:="9871";
                when 9872 => b:="9872";
                when 9873 => b:="9873";
                when 9874 => b:="9874";
                when 9875 => b:="9875";
                when 9876 => b:="9876";
                when 9877 => b:="9877";
                when 9878 => b:="9878";
                when 9879 => b:="9879";
                when 9880 => b:="9880";
                when 9881 => b:="9881";
                when 9882 => b:="9882";
                when 9883 => b:="9883";
                when 9884 => b:="9884";
                when 9885 => b:="9885";
                when 9886 => b:="9886";
                when 9887 => b:="9887";
                when 9888 => b:="9888";
                when 9889 => b:="9889";
                when 9890 => b:="9890";
                when 9891 => b:="9891";
                when 9892 => b:="9892";
                when 9893 => b:="9893";
                when 9894 => b:="9894";
                when 9895 => b:="9895";
                when 9896 => b:="9896";
                when 9897 => b:="9897";
                when 9898 => b:="9898";
                when 9899 => b:="9899";
                when 9900 => b:="9900";
                when 9901 => b:="9901";
                when 9902 => b:="9902";
                when 9903 => b:="9903";
                when 9904 => b:="9904";
                when 9905 => b:="9905";
                when 9906 => b:="9906";
                when 9907 => b:="9907";
                when 9908 => b:="9908";
                when 9909 => b:="9909";
                when 9910 => b:="9910";
                when 9911 => b:="9911";
                when 9912 => b:="9912";
                when 9913 => b:="9913";
                when 9914 => b:="9914";
                when 9915 => b:="9915";
                when 9916 => b:="9916";
                when 9917 => b:="9917";
                when 9918 => b:="9918";
                when 9919 => b:="9919";
                when 9920 => b:="9920";
                when 9921 => b:="9921";
                when 9922 => b:="9922";
                when 9923 => b:="9923";
                when 9924 => b:="9924";
                when 9925 => b:="9925";
                when 9926 => b:="9926";
                when 9927 => b:="9927";
                when 9928 => b:="9928";
                when 9929 => b:="9929";
                when 9930 => b:="9930";
                when 9931 => b:="9931";
                when 9932 => b:="9932";
                when 9933 => b:="9933";
                when 9934 => b:="9934";
                when 9935 => b:="9935";
                when 9936 => b:="9936";
                when 9937 => b:="9937";
                when 9938 => b:="9938";
                when 9939 => b:="9939";
                when 9940 => b:="9940";
                when 9941 => b:="9941";
                when 9942 => b:="9942";
                when 9943 => b:="9943";
                when 9944 => b:="9944";
                when 9945 => b:="9945";
                when 9946 => b:="9946";
                when 9947 => b:="9947";
                when 9948 => b:="9948";
                when 9949 => b:="9949";
                when 9950 => b:="9950";
                when 9951 => b:="9951";
                when 9952 => b:="9952";
                when 9953 => b:="9953";
                when 9954 => b:="9954";
                when 9955 => b:="9955";
                when 9956 => b:="9956";
                when 9957 => b:="9957";
                when 9958 => b:="9958";
                when 9959 => b:="9959";
                when 9960 => b:="9960";
                when 9961 => b:="9961";
                when 9962 => b:="9962";
                when 9963 => b:="9963";
                when 9964 => b:="9964";
                when 9965 => b:="9965";
                when 9966 => b:="9966";
                when 9967 => b:="9967";
                when 9968 => b:="9968";
                when 9969 => b:="9969";
                when 9970 => b:="9970";
                when 9971 => b:="9971";
                when 9972 => b:="9972";
                when 9973 => b:="9973";
                when 9974 => b:="9974";
                when 9975 => b:="9975";
                when 9976 => b:="9976";
                when 9977 => b:="9977";
                when 9978 => b:="9978";
                when 9979 => b:="9979";
                when 9980 => b:="9980";
                when 9981 => b:="9981";
                when 9982 => b:="9982";
                when 9983 => b:="9983";
                when 9984 => b:="9984";
                when 9985 => b:="9985";
                when 9986 => b:="9986";
                when 9987 => b:="9987";
                when 9988 => b:="9988";
                when 9989 => b:="9989";
                when 9990 => b:="9990";
                when 9991 => b:="9991";
                when 9992 => b:="9992";
                when 9993 => b:="9993";
                when 9994 => b:="9994";
                when 9995 => b:="9995";
                when 9996 => b:="9996";
                when 9997 => b:="9997";
                when 9998 => b:="9998";
                when 9999 => b:="9999";
                when others => b:= "    ";
            end case;
            return b;
    end function inttostring; -- 4 decimal
end ConverterFunctions;
